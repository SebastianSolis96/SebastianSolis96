<svg width="1376" height="476" viewBox="0 0 1376 476" fill="none" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink">
<g clip-path="url(#clip0_367_2)">
<rect width="1376" height="476" rx="20" fill="#3F3F3F"/>
<g filter="url(#filter0_b_367_2)">
<rect width="1376" height="476" fill="url(#paint0_linear_367_2)"/>
<rect x="86" y="35" width="380" height="380" fill="url(#pattern0)"/>
<path d="M564.837 127.993C564.837 126.997 564.69 126.104 564.397 125.312C564.104 124.492 563.562 123.73 562.771 123.027C561.98 122.324 560.838 121.621 559.344 120.918C557.879 120.186 555.945 119.424 553.543 118.633C550.73 117.695 548.021 116.641 545.413 115.469C542.806 114.268 540.477 112.876 538.426 111.294C536.375 109.683 534.749 107.808 533.548 105.669C532.347 103.501 531.746 100.981 531.746 98.1104C531.746 95.3564 532.361 92.8809 533.592 90.6836C534.822 88.457 536.536 86.5674 538.733 85.0146C540.96 83.4326 543.567 82.2314 546.556 81.4111C549.544 80.5615 552.811 80.1367 556.355 80.1367C561.043 80.1367 565.174 80.957 568.748 82.5977C572.352 84.209 575.164 86.5088 577.186 89.4971C579.236 92.4561 580.262 95.957 580.262 100H564.925C564.925 98.3887 564.588 96.9678 563.914 95.7373C563.27 94.5068 562.288 93.54 560.97 92.8369C559.651 92.1338 557.996 91.7822 556.004 91.7822C554.07 91.7822 552.444 92.0752 551.126 92.6611C549.808 93.2471 548.812 94.0381 548.138 95.0342C547.464 96.001 547.127 97.0703 547.127 98.2422C547.127 99.209 547.391 100.088 547.918 100.879C548.475 101.641 549.251 102.358 550.247 103.032C551.272 103.706 552.503 104.351 553.938 104.966C555.403 105.581 557.044 106.182 558.86 106.768C562.259 107.852 565.276 109.067 567.913 110.415C570.579 111.733 572.82 113.242 574.637 114.941C576.482 116.611 577.874 118.516 578.812 120.654C579.778 122.793 580.262 125.21 580.262 127.905C580.262 130.776 579.705 133.325 578.592 135.552C577.479 137.778 575.882 139.668 573.802 141.221C571.722 142.744 569.231 143.901 566.331 144.692C563.431 145.483 560.193 145.879 556.619 145.879C553.338 145.879 550.101 145.469 546.907 144.648C543.743 143.799 540.872 142.51 538.294 140.781C535.716 139.023 533.65 136.782 532.098 134.058C530.574 131.304 529.812 128.037 529.812 124.258H545.281C545.281 126.133 545.53 127.715 546.028 129.004C546.526 130.293 547.259 131.333 548.226 132.124C549.192 132.886 550.379 133.442 551.785 133.794C553.191 134.116 554.803 134.277 556.619 134.277C558.582 134.277 560.164 133.999 561.365 133.442C562.566 132.856 563.445 132.095 564.002 131.157C564.559 130.19 564.837 129.136 564.837 127.993ZM632.249 133.135V145H598.147V133.135H632.249ZM603.641 81.0156V145H588.216V81.0156H603.641ZM627.854 106.416V117.886H598.147V106.416H627.854ZM632.381 81.0156V92.9248H598.147V81.0156H632.381ZM664.681 117.798H648.201L648.113 107.69H661.473C663.875 107.69 665.794 107.427 667.229 106.899C668.665 106.343 669.705 105.537 670.35 104.482C671.023 103.428 671.36 102.109 671.36 100.527C671.36 98.7109 671.023 97.2461 670.35 96.1328C669.676 95.0195 668.606 94.2139 667.142 93.7158C665.706 93.1885 663.846 92.9248 661.561 92.9248H654.002V145H638.577V81.0156H661.561C665.516 81.0156 669.046 81.3818 672.151 82.1143C675.257 82.8174 677.894 83.9014 680.062 85.3662C682.259 86.8311 683.929 88.6768 685.071 90.9033C686.214 93.1006 686.785 95.6934 686.785 98.6816C686.785 101.289 686.229 103.735 685.115 106.021C684.002 108.306 682.142 110.166 679.534 111.602C676.956 113.008 673.426 113.74 668.943 113.799L664.681 117.798ZM664.065 145H644.466L649.739 133.135H664.065C666.175 133.135 667.859 132.812 669.119 132.168C670.408 131.494 671.331 130.615 671.888 129.531C672.474 128.418 672.767 127.188 672.767 125.84C672.767 124.199 672.488 122.778 671.932 121.577C671.404 120.376 670.555 119.453 669.383 118.809C668.211 118.135 666.644 117.798 664.681 117.798H651.717L651.805 107.69H667.317L670.921 111.733C675.198 111.558 678.582 112.158 681.072 113.535C683.592 114.912 685.394 116.729 686.478 118.984C687.562 121.24 688.104 123.599 688.104 126.06C688.104 130.249 687.195 133.75 685.379 136.562C683.592 139.375 680.911 141.484 677.337 142.891C673.763 144.297 669.339 145 664.065 145ZM723.787 94.4629L708.187 145H691.619L715.13 81.0156H725.633L723.787 94.4629ZM736.707 145L721.062 94.4629L719.041 81.0156H729.676L753.318 145H736.707ZM736.092 121.138V133.047H703.265V121.138H736.092ZM790.979 127.993C790.979 126.997 790.833 126.104 790.54 125.312C790.247 124.492 789.705 123.73 788.914 123.027C788.123 122.324 786.98 121.621 785.486 120.918C784.021 120.186 782.088 119.424 779.686 118.633C776.873 117.695 774.163 116.641 771.556 115.469C768.948 114.268 766.619 112.876 764.568 111.294C762.518 109.683 760.892 107.808 759.69 105.669C758.489 103.501 757.889 100.981 757.889 98.1104C757.889 95.3564 758.504 92.8809 759.734 90.6836C760.965 88.457 762.679 86.5674 764.876 85.0146C767.103 83.4326 769.71 82.2314 772.698 81.4111C775.687 80.5615 778.953 80.1367 782.498 80.1367C787.186 80.1367 791.316 80.957 794.891 82.5977C798.494 84.209 801.307 86.5088 803.328 89.4971C805.379 92.4561 806.404 95.957 806.404 100H791.067C791.067 98.3887 790.73 96.9678 790.057 95.7373C789.412 94.5068 788.431 93.54 787.112 92.8369C785.794 92.1338 784.139 91.7822 782.146 91.7822C780.213 91.7822 778.587 92.0752 777.269 92.6611C775.95 93.2471 774.954 94.0381 774.28 95.0342C773.606 96.001 773.27 97.0703 773.27 98.2422C773.27 99.209 773.533 100.088 774.061 100.879C774.617 101.641 775.394 102.358 776.39 103.032C777.415 103.706 778.646 104.351 780.081 104.966C781.546 105.581 783.187 106.182 785.003 106.768C788.401 107.852 791.419 109.067 794.056 110.415C796.722 111.733 798.963 113.242 800.779 114.941C802.625 116.611 804.017 118.516 804.954 120.654C805.921 122.793 806.404 125.21 806.404 127.905C806.404 130.776 805.848 133.325 804.734 135.552C803.621 137.778 802.024 139.668 799.944 141.221C797.864 142.744 795.374 143.901 792.474 144.692C789.573 145.483 786.336 145.879 782.762 145.879C779.48 145.879 776.243 145.469 773.05 144.648C769.886 143.799 767.015 142.51 764.437 140.781C761.858 139.023 759.793 136.782 758.24 134.058C756.717 131.304 755.955 128.037 755.955 124.258H771.424C771.424 126.133 771.673 127.715 772.171 129.004C772.669 130.293 773.401 131.333 774.368 132.124C775.335 132.886 776.521 133.442 777.928 133.794C779.334 134.116 780.945 134.277 782.762 134.277C784.725 134.277 786.307 133.999 787.508 133.442C788.709 132.856 789.588 132.095 790.145 131.157C790.701 130.19 790.979 129.136 790.979 127.993ZM845.34 81.0156V145H829.915V81.0156H845.34ZM864.588 81.0156V92.9248H811.106V81.0156H864.588ZM887.527 81.0156V145H872.146V81.0156H887.527ZM926.287 94.4629L910.687 145H894.119L917.63 81.0156H928.133L926.287 94.4629ZM939.207 145L923.562 94.4629L921.541 81.0156H932.176L955.818 145H939.207ZM938.592 121.138V133.047H905.765V121.138H938.592ZM1013.96 81.0156V145H998.577L975.945 105.186V145H960.521V81.0156H975.945L998.577 120.83V81.0156H1013.96ZM1079.08 127.993C1079.08 126.997 1078.94 126.104 1078.65 125.312C1078.35 124.492 1077.81 123.73 1077.02 123.027C1076.23 122.324 1075.09 121.621 1073.59 120.918C1072.13 120.186 1070.19 119.424 1067.79 118.633C1064.98 117.695 1062.27 116.641 1059.66 115.469C1057.05 114.268 1054.72 112.876 1052.67 111.294C1050.62 109.683 1049 107.808 1047.8 105.669C1046.59 103.501 1045.99 100.981 1045.99 98.1104C1045.99 95.3564 1046.61 92.8809 1047.84 90.6836C1049.07 88.457 1050.78 86.5674 1052.98 85.0146C1055.21 83.4326 1057.82 82.2314 1060.8 81.4111C1063.79 80.5615 1067.06 80.1367 1070.6 80.1367C1075.29 80.1367 1079.42 80.957 1083 82.5977C1086.6 84.209 1089.41 86.5088 1091.43 89.4971C1093.48 92.4561 1094.51 95.957 1094.51 100H1079.17C1079.17 98.3887 1078.84 96.9678 1078.16 95.7373C1077.52 94.5068 1076.54 93.54 1075.22 92.8369C1073.9 92.1338 1072.24 91.7822 1070.25 91.7822C1068.32 91.7822 1066.69 92.0752 1065.37 92.6611C1064.06 93.2471 1063.06 94.0381 1062.39 95.0342C1061.71 96.001 1061.38 97.0703 1061.38 98.2422C1061.38 99.209 1061.64 100.088 1062.17 100.879C1062.72 101.641 1063.5 102.358 1064.5 103.032C1065.52 103.706 1066.75 104.351 1068.19 104.966C1069.65 105.581 1071.29 106.182 1073.11 106.768C1076.51 107.852 1079.52 109.067 1082.16 110.415C1084.83 111.733 1087.07 113.242 1088.88 114.941C1090.73 116.611 1092.12 118.516 1093.06 120.654C1094.03 122.793 1094.51 125.21 1094.51 127.905C1094.51 130.776 1093.95 133.325 1092.84 135.552C1091.73 137.778 1090.13 139.668 1088.05 141.221C1085.97 142.744 1083.48 143.901 1080.58 144.692C1077.68 145.483 1074.44 145.879 1070.87 145.879C1067.59 145.879 1064.35 145.469 1061.16 144.648C1057.99 143.799 1055.12 142.51 1052.54 140.781C1049.96 139.023 1047.9 136.782 1046.35 134.058C1044.82 131.304 1044.06 128.037 1044.06 124.258H1059.53C1059.53 126.133 1059.78 127.715 1060.28 129.004C1060.77 130.293 1061.51 131.333 1062.47 132.124C1063.44 132.886 1064.63 133.442 1066.03 133.794C1067.44 134.116 1069.05 134.277 1070.87 134.277C1072.83 134.277 1074.41 133.999 1075.61 133.442C1076.81 132.856 1077.69 132.095 1078.25 131.157C1078.81 130.19 1079.08 129.136 1079.08 127.993ZM1156.6 111.733V114.326C1156.6 119.219 1155.92 123.613 1154.54 127.51C1153.19 131.377 1151.27 134.688 1148.78 137.441C1146.29 140.166 1143.35 142.261 1139.95 143.726C1136.55 145.161 1132.8 145.879 1128.7 145.879C1124.57 145.879 1120.79 145.161 1117.36 143.726C1113.96 142.261 1111 140.166 1108.48 137.441C1105.99 134.688 1104.06 131.377 1102.68 127.51C1101.34 123.613 1100.66 119.219 1100.66 114.326V111.733C1100.66 106.841 1101.34 102.446 1102.68 98.5498C1104.06 94.6533 1105.98 91.3428 1108.44 88.6182C1110.93 85.8643 1113.88 83.7695 1117.27 82.334C1120.7 80.8691 1124.48 80.1367 1128.61 80.1367C1132.71 80.1367 1136.46 80.8691 1139.86 82.334C1143.29 83.7695 1146.25 85.8643 1148.74 88.6182C1151.23 91.3428 1153.16 94.6533 1154.54 98.5498C1155.92 102.446 1156.6 106.841 1156.6 111.733ZM1140.96 114.326V111.646C1140.96 108.481 1140.68 105.698 1140.12 103.296C1139.6 100.864 1138.81 98.8281 1137.75 97.1875C1136.7 95.5469 1135.39 94.3164 1133.84 93.4961C1132.32 92.6465 1130.57 92.2217 1128.61 92.2217C1126.56 92.2217 1124.77 92.6465 1123.25 93.4961C1121.73 94.3164 1120.45 95.5469 1119.43 97.1875C1118.4 98.8281 1117.62 100.864 1117.1 103.296C1116.6 105.698 1116.35 108.481 1116.35 111.646V114.326C1116.35 117.461 1116.6 120.244 1117.1 122.676C1117.62 125.078 1118.4 127.114 1119.43 128.784C1120.48 130.454 1121.77 131.714 1123.29 132.563C1124.85 133.413 1126.65 133.838 1128.7 133.838C1130.66 133.838 1132.41 133.413 1133.93 132.563C1135.45 131.714 1136.73 130.454 1137.75 128.784C1138.81 127.114 1139.6 125.078 1140.12 122.676C1140.68 120.244 1140.96 117.461 1140.96 114.326ZM1206.88 133.135V145H1174.53V133.135H1206.88ZM1180.03 81.0156V145H1164.6V81.0156H1180.03ZM1229.77 81.0156V145H1214.39V81.0156H1229.77ZM1273.59 127.993C1273.59 126.997 1273.44 126.104 1273.15 125.312C1272.85 124.492 1272.31 123.73 1271.52 123.027C1270.73 122.324 1269.59 121.621 1268.09 120.918C1266.63 120.186 1264.7 119.424 1262.29 118.633C1259.48 117.695 1256.77 116.641 1254.16 115.469C1251.56 114.268 1249.23 112.876 1247.18 111.294C1245.12 109.683 1243.5 107.808 1242.3 105.669C1241.1 103.501 1240.5 100.981 1240.5 98.1104C1240.5 95.3564 1241.11 92.8809 1242.34 90.6836C1243.57 88.457 1245.29 86.5674 1247.48 85.0146C1249.71 83.4326 1252.32 82.2314 1255.31 81.4111C1258.29 80.5615 1261.56 80.1367 1265.11 80.1367C1269.79 80.1367 1273.92 80.957 1277.5 82.5977C1281.1 84.209 1283.91 86.5088 1285.94 89.4971C1287.99 92.4561 1289.01 95.957 1289.01 100H1273.67C1273.67 98.3887 1273.34 96.9678 1272.66 95.7373C1272.02 94.5068 1271.04 93.54 1269.72 92.8369C1268.4 92.1338 1266.75 91.7822 1264.75 91.7822C1262.82 91.7822 1261.19 92.0752 1259.88 92.6611C1258.56 93.2471 1257.56 94.0381 1256.89 95.0342C1256.21 96.001 1255.88 97.0703 1255.88 98.2422C1255.88 99.209 1256.14 100.088 1256.67 100.879C1257.22 101.641 1258 102.358 1259 103.032C1260.02 103.706 1261.25 104.351 1262.69 104.966C1264.15 105.581 1265.79 106.182 1267.61 106.768C1271.01 107.852 1274.03 109.067 1276.66 110.415C1279.33 111.733 1281.57 113.242 1283.39 114.941C1285.23 116.611 1286.62 118.516 1287.56 120.654C1288.53 122.793 1289.01 125.21 1289.01 127.905C1289.01 130.776 1288.46 133.325 1287.34 135.552C1286.23 137.778 1284.63 139.668 1282.55 141.221C1280.47 142.744 1277.98 143.901 1275.08 144.692C1272.18 145.483 1268.94 145.879 1265.37 145.879C1262.09 145.879 1258.85 145.469 1255.66 144.648C1252.49 143.799 1249.62 142.51 1247.04 140.781C1244.47 139.023 1242.4 136.782 1240.85 134.058C1239.32 131.304 1238.56 128.037 1238.56 124.258H1254.03C1254.03 126.133 1254.28 127.715 1254.78 129.004C1255.28 130.293 1256.01 131.333 1256.98 132.124C1257.94 132.886 1259.13 133.442 1260.54 133.794C1261.94 134.116 1263.55 134.277 1265.37 134.277C1267.33 134.277 1268.91 133.999 1270.12 133.442C1271.32 132.856 1272.2 132.095 1272.75 131.157C1273.31 130.19 1273.59 129.136 1273.59 127.993Z" fill="white"/>
<path d="M720.539 224.453V260H713.825V224.453H720.539ZM734.87 239.81V245.107H718.781V239.81H734.87ZM736.75 224.453V229.751H718.781V224.453H736.75ZM749.138 238.979V260H742.692V233.584H748.796L749.138 238.979ZM757.17 233.413L757.072 239.419C756.714 239.354 756.307 239.305 755.852 239.272C755.412 239.24 754.997 239.224 754.606 239.224C753.614 239.224 752.743 239.362 751.994 239.639C751.245 239.899 750.619 240.282 750.114 240.786C749.626 241.291 749.252 241.909 748.991 242.642C748.731 243.358 748.584 244.172 748.552 245.083L747.16 244.912C747.16 243.236 747.331 241.681 747.673 240.249C748.015 238.817 748.511 237.563 749.162 236.489C749.813 235.415 750.627 234.585 751.604 233.999C752.596 233.397 753.736 233.096 755.021 233.096C755.38 233.096 755.762 233.128 756.169 233.193C756.592 233.242 756.926 233.315 757.17 233.413ZM761.379 247.061V246.548C761.379 244.611 761.656 242.829 762.209 241.201C762.762 239.557 763.568 238.133 764.626 236.929C765.684 235.724 766.978 234.788 768.508 234.121C770.038 233.438 771.779 233.096 773.732 233.096C775.718 233.096 777.476 233.438 779.006 234.121C780.552 234.788 781.854 235.724 782.912 236.929C783.97 238.133 784.776 239.557 785.329 241.201C785.882 242.829 786.159 244.611 786.159 246.548V247.061C786.159 248.981 785.882 250.763 785.329 252.407C784.776 254.035 783.97 255.459 782.912 256.68C781.854 257.884 780.56 258.82 779.03 259.487C777.5 260.155 775.751 260.488 773.781 260.488C771.828 260.488 770.078 260.155 768.532 259.487C766.986 258.82 765.684 257.884 764.626 256.68C763.568 255.459 762.762 254.035 762.209 252.407C761.656 250.763 761.379 248.981 761.379 247.061ZM767.824 246.548V247.061C767.824 248.216 767.938 249.299 768.166 250.308C768.394 251.317 768.744 252.204 769.216 252.969C769.688 253.734 770.298 254.336 771.047 254.775C771.812 255.199 772.723 255.41 773.781 255.41C774.823 255.41 775.718 255.199 776.467 254.775C777.215 254.336 777.826 253.734 778.298 252.969C778.786 252.204 779.144 251.317 779.372 250.308C779.6 249.299 779.714 248.216 779.714 247.061V246.548C779.714 245.409 779.6 244.342 779.372 243.35C779.144 242.34 778.786 241.453 778.298 240.688C777.826 239.907 777.207 239.297 776.442 238.857C775.694 238.402 774.79 238.174 773.732 238.174C772.691 238.174 771.796 238.402 771.047 238.857C770.298 239.297 769.688 239.907 769.216 240.688C768.744 241.453 768.394 242.34 768.166 243.35C767.938 244.342 767.824 245.409 767.824 246.548ZM799.67 239.224V260H793.225V233.584H799.279L799.67 239.224ZM798.645 245.84H796.74C796.757 243.919 797.017 242.178 797.521 240.615C798.026 239.053 798.734 237.71 799.646 236.587C800.573 235.464 801.672 234.601 802.941 233.999C804.211 233.397 805.627 233.096 807.189 233.096C808.459 233.096 809.606 233.275 810.632 233.633C811.657 233.991 812.536 234.561 813.269 235.342C814.017 236.123 814.587 237.148 814.978 238.418C815.384 239.671 815.588 241.217 815.588 243.057V260H809.094V243.008C809.094 241.803 808.915 240.851 808.557 240.151C808.215 239.451 807.71 238.955 807.043 238.662C806.392 238.369 805.586 238.223 804.626 238.223C803.633 238.223 802.762 238.426 802.014 238.833C801.281 239.224 800.663 239.769 800.158 240.469C799.67 241.169 799.296 241.974 799.035 242.886C798.775 243.797 798.645 244.782 798.645 245.84ZM836.276 233.584V238.223H821.14V233.584H836.276ZM825.192 227.09H831.662V252.383C831.662 253.164 831.768 253.766 831.979 254.189C832.191 254.613 832.508 254.897 832.932 255.044C833.355 255.19 833.859 255.264 834.445 255.264C834.868 255.264 835.259 255.239 835.617 255.19C835.975 255.142 836.276 255.093 836.521 255.044L836.545 259.878C836.008 260.057 835.397 260.203 834.714 260.317C834.047 260.431 833.29 260.488 832.443 260.488C830.995 260.488 829.725 260.244 828.635 259.756C827.544 259.251 826.698 258.446 826.096 257.339C825.493 256.216 825.192 254.735 825.192 252.896V227.09ZM854.938 260.488C852.937 260.488 851.138 260.163 849.543 259.512C847.948 258.861 846.589 257.957 845.466 256.802C844.359 255.63 843.505 254.271 842.902 252.725C842.316 251.162 842.023 249.486 842.023 247.695V246.719C842.023 244.684 842.316 242.837 842.902 241.177C843.488 239.5 844.318 238.06 845.393 236.855C846.467 235.651 847.753 234.723 849.25 234.072C850.747 233.421 852.399 233.096 854.206 233.096C856.078 233.096 857.73 233.413 859.162 234.048C860.594 234.666 861.791 235.545 862.751 236.685C863.711 237.824 864.436 239.191 864.924 240.786C865.412 242.365 865.656 244.115 865.656 246.035V248.745H844.953V244.302H859.309V243.813C859.276 242.788 859.081 241.852 858.723 241.006C858.365 240.143 857.811 239.46 857.062 238.955C856.314 238.434 855.345 238.174 854.157 238.174C853.197 238.174 852.359 238.385 851.643 238.809C850.943 239.215 850.357 239.801 849.885 240.566C849.429 241.315 849.087 242.21 848.859 243.252C848.632 244.294 848.518 245.449 848.518 246.719V247.695C848.518 248.802 848.664 249.827 848.957 250.771C849.266 251.715 849.714 252.537 850.3 253.237C850.902 253.921 851.618 254.458 852.448 254.849C853.295 255.223 854.255 255.41 855.329 255.41C856.68 255.41 857.901 255.15 858.991 254.629C860.098 254.092 861.058 253.302 861.872 252.261L865.119 255.63C864.566 256.444 863.817 257.225 862.873 257.974C861.945 258.722 860.822 259.333 859.504 259.805C858.186 260.26 856.664 260.488 854.938 260.488ZM878.801 239.224V260H872.355V233.584H878.41L878.801 239.224ZM877.775 245.84H875.871C875.887 243.919 876.148 242.178 876.652 240.615C877.157 239.053 877.865 237.71 878.776 236.587C879.704 235.464 880.803 234.601 882.072 233.999C883.342 233.397 884.758 233.096 886.32 233.096C887.59 233.096 888.737 233.275 889.763 233.633C890.788 233.991 891.667 234.561 892.399 235.342C893.148 236.123 893.718 237.148 894.108 238.418C894.515 239.671 894.719 241.217 894.719 243.057V260H888.225V243.008C888.225 241.803 888.046 240.851 887.688 240.151C887.346 239.451 886.841 238.955 886.174 238.662C885.523 238.369 884.717 238.223 883.757 238.223C882.764 238.223 881.893 238.426 881.145 238.833C880.412 239.224 879.794 239.769 879.289 240.469C878.801 241.169 878.426 241.974 878.166 242.886C877.906 243.797 877.775 244.782 877.775 245.84ZM918.752 254.385V222.5H925.246V260H919.387L918.752 254.385ZM901.784 247.109V246.597C901.784 244.578 902.012 242.747 902.468 241.104C902.94 239.443 903.623 238.019 904.519 236.831C905.414 235.643 906.496 234.723 907.766 234.072C909.051 233.421 910.508 233.096 912.136 233.096C913.715 233.096 915.09 233.413 916.262 234.048C917.45 234.683 918.459 235.586 919.289 236.758C920.135 237.93 920.811 239.321 921.315 240.933C921.82 242.528 922.186 244.285 922.414 246.206V247.598C922.186 249.469 921.82 251.187 921.315 252.749C920.811 254.312 920.135 255.679 919.289 256.851C918.459 258.006 917.45 258.901 916.262 259.536C915.074 260.171 913.682 260.488 912.087 260.488C910.476 260.488 909.027 260.155 907.741 259.487C906.472 258.82 905.389 257.884 904.494 256.68C903.615 255.475 902.94 254.059 902.468 252.432C902.012 250.804 901.784 249.03 901.784 247.109ZM908.254 246.597V247.109C908.254 248.249 908.352 249.315 908.547 250.308C908.742 251.3 909.06 252.179 909.499 252.944C909.938 253.693 910.5 254.279 911.184 254.702C911.883 255.125 912.73 255.337 913.723 255.337C914.992 255.337 916.034 255.06 916.848 254.507C917.678 253.937 918.321 253.164 918.776 252.188C919.232 251.195 919.525 250.08 919.655 248.843V245.01C919.59 244.033 919.419 243.13 919.143 242.3C918.882 241.47 918.508 240.754 918.02 240.151C917.548 239.549 916.962 239.077 916.262 238.735C915.562 238.394 914.732 238.223 913.771 238.223C912.779 238.223 911.932 238.442 911.232 238.882C910.533 239.305 909.963 239.899 909.523 240.664C909.084 241.429 908.758 242.316 908.547 243.325C908.352 244.334 908.254 245.425 908.254 246.597ZM959.641 260H951.975L952.023 254.727H959.641C961.708 254.727 963.441 254.271 964.841 253.359C966.241 252.432 967.299 251.105 968.015 249.38C968.731 247.638 969.089 245.555 969.089 243.13V241.299C969.089 239.427 968.885 237.775 968.479 236.343C968.072 234.91 967.469 233.706 966.672 232.729C965.891 231.753 964.922 231.012 963.767 230.508C962.611 230.003 961.285 229.751 959.787 229.751H951.828V224.453H959.787C962.163 224.453 964.328 224.852 966.281 225.649C968.251 226.447 969.951 227.594 971.384 229.092C972.832 230.573 973.939 232.347 974.704 234.414C975.485 236.481 975.876 238.792 975.876 241.348V243.13C975.876 245.669 975.485 247.98 974.704 250.063C973.939 252.131 972.832 253.905 971.384 255.386C969.951 256.867 968.243 258.006 966.257 258.804C964.271 259.601 962.066 260 959.641 260ZM955.734 224.453V260H949.021V224.453H955.734ZM995.466 260.488C993.464 260.488 991.665 260.163 990.07 259.512C988.475 258.861 987.116 257.957 985.993 256.802C984.886 255.63 984.032 254.271 983.43 252.725C982.844 251.162 982.551 249.486 982.551 247.695V246.719C982.551 244.684 982.844 242.837 983.43 241.177C984.016 239.5 984.846 238.06 985.92 236.855C986.994 235.651 988.28 234.723 989.777 234.072C991.275 233.421 992.927 233.096 994.733 233.096C996.605 233.096 998.257 233.413 999.689 234.048C1001.12 234.666 1002.32 235.545 1003.28 236.685C1004.24 237.824 1004.96 239.191 1005.45 240.786C1005.94 242.365 1006.18 244.115 1006.18 246.035V248.745H985.48V244.302H999.836V243.813C999.803 242.788 999.608 241.852 999.25 241.006C998.892 240.143 998.339 239.46 997.59 238.955C996.841 238.434 995.873 238.174 994.685 238.174C993.724 238.174 992.886 238.385 992.17 238.809C991.47 239.215 990.884 239.801 990.412 240.566C989.956 241.315 989.615 242.21 989.387 243.252C989.159 244.294 989.045 245.449 989.045 246.719V247.695C989.045 248.802 989.191 249.827 989.484 250.771C989.794 251.715 990.241 252.537 990.827 253.237C991.429 253.921 992.146 254.458 992.976 254.849C993.822 255.223 994.782 255.41 995.856 255.41C997.207 255.41 998.428 255.15 999.519 254.629C1000.63 254.092 1001.59 253.302 1002.4 252.261L1005.65 255.63C1005.09 256.444 1004.34 257.225 1003.4 257.974C1002.47 258.722 1001.35 259.333 1000.03 259.805C998.713 260.26 997.191 260.488 995.466 260.488ZM1021.43 255.117L1027.58 233.584H1034.32L1025.26 260H1021.16L1021.43 255.117ZM1016.94 233.584L1023.16 255.166L1023.38 260H1019.25L1010.17 233.584H1016.94ZM1051.74 260.488C1049.73 260.488 1047.93 260.163 1046.34 259.512C1044.74 258.861 1043.39 257.957 1042.26 256.802C1041.16 255.63 1040.3 254.271 1039.7 252.725C1039.11 251.162 1038.82 249.486 1038.82 247.695V246.719C1038.82 244.684 1039.11 242.837 1039.7 241.177C1040.29 239.5 1041.12 238.06 1042.19 236.855C1043.26 235.651 1044.55 234.723 1046.05 234.072C1047.54 233.421 1049.2 233.096 1051 233.096C1052.87 233.096 1054.53 233.413 1055.96 234.048C1057.39 234.666 1058.59 235.545 1059.55 236.685C1060.51 237.824 1061.23 239.191 1061.72 240.786C1062.21 242.365 1062.45 244.115 1062.45 246.035V248.745H1041.75V244.302H1056.11V243.813C1056.07 242.788 1055.88 241.852 1055.52 241.006C1055.16 240.143 1054.61 239.46 1053.86 238.955C1053.11 238.434 1052.14 238.174 1050.95 238.174C1049.99 238.174 1049.16 238.385 1048.44 238.809C1047.74 239.215 1047.15 239.801 1046.68 240.566C1046.23 241.315 1045.88 242.21 1045.66 243.252C1045.43 244.294 1045.31 245.449 1045.31 246.719V247.695C1045.31 248.802 1045.46 249.827 1045.75 250.771C1046.06 251.715 1046.51 252.537 1047.1 253.237C1047.7 253.921 1048.42 254.458 1049.25 254.849C1050.09 255.223 1051.05 255.41 1052.13 255.41C1053.48 255.41 1054.7 255.15 1055.79 254.629C1056.89 254.092 1057.86 253.302 1058.67 252.261L1061.92 255.63C1061.36 256.444 1060.61 257.225 1059.67 257.974C1058.74 258.722 1057.62 259.333 1056.3 259.805C1054.98 260.26 1053.46 260.488 1051.74 260.488ZM1076.11 222.5V260H1069.64V222.5H1076.11ZM1083.62 247.061V246.548C1083.62 244.611 1083.89 242.829 1084.45 241.201C1085 239.557 1085.8 238.133 1086.86 236.929C1087.92 235.724 1089.21 234.788 1090.74 234.121C1092.27 233.438 1094.02 233.096 1095.97 233.096C1097.95 233.096 1099.71 233.438 1101.24 234.121C1102.79 234.788 1104.09 235.724 1105.15 236.929C1106.21 238.133 1107.01 239.557 1107.57 241.201C1108.12 242.829 1108.4 244.611 1108.4 246.548V247.061C1108.4 248.981 1108.12 250.763 1107.57 252.407C1107.01 254.035 1106.21 255.459 1105.15 256.68C1104.09 257.884 1102.8 258.82 1101.27 259.487C1099.74 260.155 1097.99 260.488 1096.02 260.488C1094.06 260.488 1092.31 260.155 1090.77 259.487C1089.22 258.82 1087.92 257.884 1086.86 256.68C1085.8 255.459 1085 254.035 1084.45 252.407C1083.89 250.763 1083.62 248.981 1083.62 247.061ZM1090.06 246.548V247.061C1090.06 248.216 1090.17 249.299 1090.4 250.308C1090.63 251.317 1090.98 252.204 1091.45 252.969C1091.92 253.734 1092.53 254.336 1093.28 254.775C1094.05 255.199 1094.96 255.41 1096.02 255.41C1097.06 255.41 1097.95 255.199 1098.7 254.775C1099.45 254.336 1100.06 253.734 1100.53 252.969C1101.02 252.204 1101.38 251.317 1101.61 250.308C1101.84 249.299 1101.95 248.216 1101.95 247.061V246.548C1101.95 245.409 1101.84 244.342 1101.61 243.35C1101.38 242.34 1101.02 241.453 1100.53 240.688C1100.06 239.907 1099.44 239.297 1098.68 238.857C1097.93 238.402 1097.03 238.174 1095.97 238.174C1094.93 238.174 1094.03 238.402 1093.28 238.857C1092.53 239.297 1091.92 239.907 1091.45 240.688C1090.98 241.453 1090.63 242.34 1090.4 243.35C1090.17 244.342 1090.06 245.409 1090.06 246.548ZM1122.03 238.662V270.156H1115.56V233.584H1121.54L1122.03 238.662ZM1139 246.523V247.036C1139 248.957 1138.77 250.739 1138.31 252.383C1137.87 254.01 1137.22 255.435 1136.36 256.655C1135.5 257.86 1134.42 258.804 1133.14 259.487C1131.87 260.155 1130.4 260.488 1128.74 260.488C1127.11 260.488 1125.7 260.179 1124.49 259.561C1123.29 258.926 1122.27 258.031 1121.44 256.875C1120.61 255.719 1119.94 254.377 1119.44 252.847C1118.95 251.3 1118.59 249.616 1118.34 247.793V246.157C1118.59 244.22 1118.95 242.463 1119.44 240.884C1119.94 239.289 1120.61 237.913 1121.44 236.758C1122.27 235.586 1123.28 234.683 1124.47 234.048C1125.67 233.413 1127.08 233.096 1128.69 233.096C1130.37 233.096 1131.84 233.413 1133.11 234.048C1134.4 234.683 1135.48 235.594 1136.36 236.782C1137.24 237.97 1137.9 239.386 1138.34 241.03C1138.78 242.674 1139 244.505 1139 246.523ZM1132.53 247.036V246.523C1132.53 245.352 1132.42 244.269 1132.21 243.276C1132 242.267 1131.67 241.388 1131.23 240.64C1130.79 239.875 1130.22 239.281 1129.52 238.857C1128.82 238.434 1127.98 238.223 1126.98 238.223C1125.99 238.223 1125.14 238.385 1124.42 238.711C1123.7 239.036 1123.12 239.5 1122.66 240.103C1122.21 240.705 1121.85 241.421 1121.59 242.251C1121.34 243.065 1121.18 243.968 1121.1 244.961V249.014C1121.25 250.218 1121.53 251.3 1121.96 252.261C1122.38 253.221 1123 253.986 1123.81 254.556C1124.64 255.125 1125.71 255.41 1127.03 255.41C1128.03 255.41 1128.87 255.19 1129.57 254.751C1130.27 254.312 1130.84 253.709 1131.28 252.944C1131.72 252.163 1132.04 251.268 1132.23 250.259C1132.43 249.25 1132.53 248.175 1132.53 247.036ZM1158.07 260.488C1156.07 260.488 1154.27 260.163 1152.68 259.512C1151.08 258.861 1149.72 257.957 1148.6 256.802C1147.49 255.63 1146.64 254.271 1146.04 252.725C1145.45 251.162 1145.16 249.486 1145.16 247.695V246.719C1145.16 244.684 1145.45 242.837 1146.04 241.177C1146.62 239.5 1147.45 238.06 1148.53 236.855C1149.6 235.651 1150.89 234.723 1152.38 234.072C1153.88 233.421 1155.53 233.096 1157.34 233.096C1159.21 233.096 1160.86 233.413 1162.3 234.048C1163.73 234.666 1164.93 235.545 1165.89 236.685C1166.85 237.824 1167.57 239.191 1168.06 240.786C1168.55 242.365 1168.79 244.115 1168.79 246.035V248.745H1148.09V244.302H1162.44V243.813C1162.41 242.788 1162.22 241.852 1161.86 241.006C1161.5 240.143 1160.95 239.46 1160.2 238.955C1159.45 238.434 1158.48 238.174 1157.29 238.174C1156.33 238.174 1155.49 238.385 1154.78 238.809C1154.08 239.215 1153.49 239.801 1153.02 240.566C1152.56 241.315 1152.22 242.21 1151.99 243.252C1151.77 244.294 1151.65 245.449 1151.65 246.719V247.695C1151.65 248.802 1151.8 249.827 1152.09 250.771C1152.4 251.715 1152.85 252.537 1153.43 253.237C1154.04 253.921 1154.75 254.458 1155.58 254.849C1156.43 255.223 1157.39 255.41 1158.46 255.41C1159.81 255.41 1161.04 255.15 1162.13 254.629C1163.23 254.092 1164.19 253.302 1165.01 252.261L1168.25 255.63C1167.7 256.444 1166.95 257.225 1166.01 257.974C1165.08 258.722 1163.96 259.333 1162.64 259.805C1161.32 260.26 1159.8 260.488 1158.07 260.488ZM1182.06 238.979V260H1175.61V233.584H1181.72L1182.06 238.979ZM1190.09 233.413L1189.99 239.419C1189.63 239.354 1189.23 239.305 1188.77 239.272C1188.33 239.24 1187.92 239.224 1187.53 239.224C1186.53 239.224 1185.66 239.362 1184.91 239.639C1184.17 239.899 1183.54 240.282 1183.03 240.786C1182.55 241.291 1182.17 241.909 1181.91 242.642C1181.65 243.358 1181.5 244.172 1181.47 245.083L1180.08 244.912C1180.08 243.236 1180.25 241.681 1180.59 240.249C1180.93 238.817 1181.43 237.563 1182.08 236.489C1182.73 235.415 1183.55 234.585 1184.52 233.999C1185.52 233.397 1186.66 233.096 1187.94 233.096C1188.3 233.096 1188.68 233.128 1189.09 233.193C1189.51 233.242 1189.85 233.315 1190.09 233.413ZM1221.92 255.41C1222.83 255.41 1223.65 255.231 1224.36 254.873C1225.08 254.515 1225.65 254.01 1226.07 253.359C1226.51 252.708 1226.75 251.951 1226.78 251.089H1232.86C1232.83 252.879 1232.32 254.482 1231.34 255.898C1230.37 257.314 1229.07 258.438 1227.44 259.268C1225.83 260.081 1224.02 260.488 1222.02 260.488C1219.98 260.488 1218.21 260.146 1216.7 259.463C1215.18 258.779 1213.92 257.827 1212.91 256.606C1211.92 255.386 1211.17 253.97 1210.67 252.358C1210.18 250.747 1209.93 249.022 1209.93 247.183V246.401C1209.93 244.562 1210.18 242.837 1210.67 241.226C1211.17 239.614 1211.92 238.198 1212.91 236.978C1213.92 235.757 1215.18 234.805 1216.7 234.121C1218.21 233.438 1219.98 233.096 1221.99 233.096C1224.13 233.096 1226 233.511 1227.61 234.341C1229.24 235.171 1230.51 236.343 1231.42 237.856C1232.35 239.37 1232.83 241.152 1232.86 243.203H1226.78C1226.75 242.259 1226.54 241.413 1226.14 240.664C1225.75 239.915 1225.2 239.313 1224.48 238.857C1223.77 238.402 1222.9 238.174 1221.87 238.174C1220.78 238.174 1219.87 238.402 1219.14 238.857C1218.42 239.313 1217.86 239.94 1217.45 240.737C1217.06 241.519 1216.79 242.397 1216.62 243.374C1216.48 244.334 1216.4 245.343 1216.4 246.401V247.183C1216.4 248.257 1216.48 249.282 1216.62 250.259C1216.79 251.235 1217.06 252.114 1217.45 252.896C1217.86 253.66 1218.42 254.271 1219.14 254.727C1219.87 255.182 1220.8 255.41 1221.92 255.41ZM1238.51 247.061V246.548C1238.51 244.611 1238.78 242.829 1239.34 241.201C1239.89 239.557 1240.7 238.133 1241.75 236.929C1242.81 235.724 1244.11 234.788 1245.64 234.121C1247.17 233.438 1248.91 233.096 1250.86 233.096C1252.85 233.096 1254.6 233.438 1256.13 234.121C1257.68 234.788 1258.98 235.724 1260.04 236.929C1261.1 238.133 1261.9 239.557 1262.46 241.201C1263.01 242.829 1263.29 244.611 1263.29 246.548V247.061C1263.29 248.981 1263.01 250.763 1262.46 252.407C1261.9 254.035 1261.1 255.459 1260.04 256.68C1258.98 257.884 1257.69 258.82 1256.16 259.487C1254.63 260.155 1252.88 260.488 1250.91 260.488C1248.96 260.488 1247.21 260.155 1245.66 259.487C1244.11 258.82 1242.81 257.884 1241.75 256.68C1240.7 255.459 1239.89 254.035 1239.34 252.407C1238.78 250.763 1238.51 248.981 1238.51 247.061ZM1244.95 246.548V247.061C1244.95 248.216 1245.07 249.299 1245.29 250.308C1245.52 251.317 1245.87 252.204 1246.34 252.969C1246.82 253.734 1247.43 254.336 1248.18 254.775C1248.94 255.199 1249.85 255.41 1250.91 255.41C1251.95 255.41 1252.85 255.199 1253.6 254.775C1254.34 254.336 1254.95 253.734 1255.43 252.969C1255.92 252.204 1256.27 251.317 1256.5 250.308C1256.73 249.299 1256.84 248.216 1256.84 247.061V246.548C1256.84 245.409 1256.73 244.342 1256.5 243.35C1256.27 242.34 1255.92 241.453 1255.43 240.688C1254.95 239.907 1254.34 239.297 1253.57 238.857C1252.82 238.402 1251.92 238.174 1250.86 238.174C1249.82 238.174 1248.92 238.402 1248.18 238.857C1247.43 239.297 1246.82 239.907 1246.34 240.688C1245.87 241.453 1245.52 242.34 1245.29 243.35C1245.07 244.342 1244.95 245.409 1244.95 246.548ZM1276.8 239.224V260H1270.35V233.584H1276.41L1276.8 239.224ZM1275.77 245.84H1273.87C1273.89 243.919 1274.15 242.178 1274.65 240.615C1275.15 239.053 1275.86 237.71 1276.77 236.587C1277.7 235.464 1278.8 234.601 1280.07 233.999C1281.34 233.397 1282.76 233.096 1284.32 233.096C1285.59 233.096 1286.74 233.275 1287.76 233.633C1288.79 233.991 1289.67 234.561 1290.4 235.342C1291.15 236.123 1291.72 237.148 1292.11 238.418C1292.51 239.671 1292.72 241.217 1292.72 243.057V260H1286.22V243.008C1286.22 241.803 1286.04 240.851 1285.69 240.151C1285.34 239.451 1284.84 238.955 1284.17 238.662C1283.52 238.369 1282.72 238.223 1281.75 238.223C1280.76 238.223 1279.89 238.426 1279.14 238.833C1278.41 239.224 1277.79 239.769 1277.29 240.469C1276.8 241.169 1276.42 241.974 1276.16 242.886C1275.9 243.797 1275.77 244.782 1275.77 245.84ZM654.47 325.41C655.381 325.41 656.195 325.231 656.911 324.873C657.627 324.515 658.197 324.01 658.62 323.359C659.06 322.708 659.296 321.951 659.328 321.089H665.407C665.375 322.879 664.87 324.482 663.894 325.898C662.917 327.314 661.615 328.438 659.987 329.268C658.376 330.081 656.569 330.488 654.567 330.488C652.533 330.488 650.759 330.146 649.245 329.463C647.731 328.779 646.47 327.827 645.461 326.606C644.468 325.386 643.719 323.97 643.215 322.358C642.727 320.747 642.482 319.022 642.482 317.183V316.401C642.482 314.562 642.727 312.837 643.215 311.226C643.719 309.614 644.468 308.198 645.461 306.978C646.47 305.757 647.731 304.805 649.245 304.121C650.759 303.438 652.525 303.096 654.543 303.096C656.675 303.096 658.547 303.511 660.158 304.341C661.786 305.171 663.055 306.343 663.967 307.856C664.895 309.37 665.375 311.152 665.407 313.203H659.328C659.296 312.259 659.084 311.413 658.693 310.664C658.303 309.915 657.749 309.313 657.033 308.857C656.317 308.402 655.446 308.174 654.421 308.174C653.33 308.174 652.419 308.402 651.687 308.857C650.97 309.313 650.409 309.94 650.002 310.737C649.611 311.519 649.335 312.397 649.172 313.374C649.025 314.334 648.952 315.343 648.952 316.401V317.183C648.952 318.257 649.025 319.282 649.172 320.259C649.335 321.235 649.611 322.114 650.002 322.896C650.409 323.66 650.97 324.271 651.687 324.727C652.419 325.182 653.347 325.41 654.47 325.41ZM687.927 323.726V303.584H694.421V330H688.317L687.927 323.726ZM688.757 318.257L690.759 318.208C690.759 319.982 690.563 321.618 690.173 323.115C689.782 324.613 689.172 325.915 688.342 327.021C687.528 328.112 686.494 328.966 685.241 329.585C683.988 330.187 682.507 330.488 680.798 330.488C679.496 330.488 678.308 330.309 677.233 329.951C676.159 329.577 675.231 328.999 674.45 328.218C673.685 327.42 673.091 326.403 672.668 325.166C672.245 323.913 672.033 322.407 672.033 320.649V303.584H678.479V320.698C678.479 321.577 678.576 322.31 678.771 322.896C678.983 323.481 679.268 323.962 679.626 324.336C680 324.694 680.432 324.954 680.92 325.117C681.424 325.264 681.962 325.337 682.531 325.337C684.094 325.337 685.323 325.028 686.218 324.409C687.129 323.774 687.78 322.928 688.171 321.87C688.562 320.796 688.757 319.591 688.757 318.257ZM709.079 308.979V330H702.634V303.584H708.737L709.079 308.979ZM717.111 303.413L717.014 309.419C716.656 309.354 716.249 309.305 715.793 309.272C715.354 309.24 714.938 309.224 714.548 309.224C713.555 309.224 712.684 309.362 711.936 309.639C711.187 309.899 710.56 310.282 710.056 310.786C709.567 311.291 709.193 311.909 708.933 312.642C708.672 313.358 708.526 314.172 708.493 315.083L707.102 314.912C707.102 313.236 707.272 311.681 707.614 310.249C707.956 308.817 708.452 307.563 709.104 306.489C709.755 305.415 710.568 304.585 711.545 303.999C712.538 303.397 713.677 303.096 714.963 303.096C715.321 303.096 715.703 303.128 716.11 303.193C716.534 303.242 716.867 303.315 717.111 303.413ZM729.987 303.584V330H723.518V303.584H729.987ZM723.078 296.675C723.078 295.715 723.404 294.917 724.055 294.282C724.722 293.647 725.617 293.33 726.74 293.33C727.863 293.33 728.75 293.647 729.401 294.282C730.069 294.917 730.402 295.715 730.402 296.675C730.402 297.619 730.069 298.408 729.401 299.043C728.75 299.678 727.863 299.995 726.74 299.995C725.617 299.995 724.722 299.678 724.055 299.043C723.404 298.408 723.078 297.619 723.078 296.675ZM737.492 317.061V316.548C737.492 314.611 737.769 312.829 738.322 311.201C738.876 309.557 739.681 308.133 740.739 306.929C741.797 305.724 743.091 304.788 744.621 304.121C746.151 303.438 747.893 303.096 749.846 303.096C751.831 303.096 753.589 303.438 755.119 304.121C756.665 304.788 757.967 305.724 759.025 306.929C760.083 308.133 760.889 309.557 761.442 311.201C761.996 312.829 762.272 314.611 762.272 316.548V317.061C762.272 318.981 761.996 320.763 761.442 322.407C760.889 324.035 760.083 325.459 759.025 326.68C757.967 327.884 756.674 328.82 755.144 329.487C753.614 330.155 751.864 330.488 749.895 330.488C747.941 330.488 746.192 330.155 744.646 329.487C743.099 328.82 741.797 327.884 740.739 326.68C739.681 325.459 738.876 324.035 738.322 322.407C737.769 320.763 737.492 318.981 737.492 317.061ZM743.938 316.548V317.061C743.938 318.216 744.051 319.299 744.279 320.308C744.507 321.317 744.857 322.204 745.329 322.969C745.801 323.734 746.411 324.336 747.16 324.775C747.925 325.199 748.837 325.41 749.895 325.41C750.936 325.41 751.831 325.199 752.58 324.775C753.329 324.336 753.939 323.734 754.411 322.969C754.899 322.204 755.257 321.317 755.485 320.308C755.713 319.299 755.827 318.216 755.827 317.061V316.548C755.827 315.409 755.713 314.342 755.485 313.35C755.257 312.34 754.899 311.453 754.411 310.688C753.939 309.907 753.321 309.297 752.556 308.857C751.807 308.402 750.904 308.174 749.846 308.174C748.804 308.174 747.909 308.402 747.16 308.857C746.411 309.297 745.801 309.907 745.329 310.688C744.857 311.453 744.507 312.34 744.279 313.35C744.051 314.342 743.938 315.409 743.938 316.548ZM783.986 322.773C783.986 322.22 783.84 321.724 783.547 321.284C783.254 320.845 782.701 320.446 781.887 320.088C781.089 319.714 779.917 319.364 778.371 319.038C777.004 318.745 775.743 318.379 774.587 317.939C773.431 317.5 772.438 316.971 771.608 316.353C770.778 315.718 770.127 314.977 769.655 314.131C769.2 313.268 768.972 312.275 768.972 311.152C768.972 310.062 769.208 309.036 769.68 308.076C770.152 307.1 770.835 306.245 771.73 305.513C772.626 304.764 773.716 304.178 775.002 303.755C776.288 303.315 777.736 303.096 779.348 303.096C781.594 303.096 783.522 303.462 785.134 304.194C786.761 304.927 788.007 305.936 788.869 307.222C789.732 308.491 790.163 309.924 790.163 311.519H783.718C783.718 310.819 783.555 310.184 783.229 309.614C782.92 309.045 782.44 308.589 781.789 308.247C781.138 307.889 780.316 307.71 779.323 307.71C778.428 307.71 777.671 307.856 777.053 308.149C776.451 308.442 775.995 308.825 775.686 309.297C775.376 309.769 775.222 310.29 775.222 310.859C775.222 311.283 775.303 311.665 775.466 312.007C775.645 312.332 775.93 312.633 776.32 312.91C776.711 313.187 777.24 313.439 777.907 313.667C778.591 313.895 779.429 314.115 780.422 314.326C782.391 314.717 784.108 315.238 785.573 315.889C787.054 316.523 788.21 317.37 789.04 318.428C789.87 319.486 790.285 320.837 790.285 322.48C790.285 323.652 790.033 324.727 789.528 325.703C789.024 326.663 788.291 327.502 787.331 328.218C786.371 328.934 785.223 329.495 783.889 329.902C782.554 330.293 781.049 330.488 779.372 330.488C776.947 330.488 774.896 330.057 773.22 329.194C771.543 328.315 770.274 327.209 769.411 325.874C768.549 324.523 768.117 323.123 768.117 321.675H774.294C774.343 322.7 774.619 323.522 775.124 324.141C775.629 324.759 776.263 325.207 777.028 325.483C777.81 325.744 778.632 325.874 779.494 325.874C780.471 325.874 781.293 325.744 781.96 325.483C782.627 325.207 783.132 324.84 783.474 324.385C783.815 323.913 783.986 323.376 783.986 322.773ZM804.528 303.584V330H798.059V303.584H804.528ZM797.619 296.675C797.619 295.715 797.945 294.917 798.596 294.282C799.263 293.647 800.158 293.33 801.281 293.33C802.404 293.33 803.291 293.647 803.942 294.282C804.61 294.917 804.943 295.715 804.943 296.675C804.943 297.619 804.61 298.408 803.942 299.043C803.291 299.678 802.404 299.995 801.281 299.995C800.158 299.995 799.263 299.678 798.596 299.043C797.945 298.408 797.619 297.619 797.619 296.675ZM829.025 324.385V292.5H835.52V330H829.66L829.025 324.385ZM812.058 317.109V316.597C812.058 314.578 812.285 312.747 812.741 311.104C813.213 309.443 813.897 308.019 814.792 306.831C815.687 305.643 816.77 304.723 818.039 304.072C819.325 303.421 820.782 303.096 822.409 303.096C823.988 303.096 825.363 303.413 826.535 304.048C827.723 304.683 828.732 305.586 829.562 306.758C830.409 307.93 831.084 309.321 831.589 310.933C832.093 312.528 832.46 314.285 832.688 316.206V317.598C832.46 319.469 832.093 321.187 831.589 322.749C831.084 324.312 830.409 325.679 829.562 326.851C828.732 328.006 827.723 328.901 826.535 329.536C825.347 330.171 823.955 330.488 822.36 330.488C820.749 330.488 819.3 330.155 818.015 329.487C816.745 328.82 815.663 327.884 814.768 326.68C813.889 325.475 813.213 324.059 812.741 322.432C812.285 320.804 812.058 319.03 812.058 317.109ZM818.527 316.597V317.109C818.527 318.249 818.625 319.315 818.82 320.308C819.016 321.3 819.333 322.179 819.772 322.944C820.212 323.693 820.773 324.279 821.457 324.702C822.157 325.125 823.003 325.337 823.996 325.337C825.266 325.337 826.307 325.06 827.121 324.507C827.951 323.937 828.594 323.164 829.05 322.188C829.506 321.195 829.799 320.08 829.929 318.843V315.01C829.864 314.033 829.693 313.13 829.416 312.3C829.156 311.47 828.781 310.754 828.293 310.151C827.821 309.549 827.235 309.077 826.535 308.735C825.835 308.394 825.005 308.223 824.045 308.223C823.052 308.223 822.206 308.442 821.506 308.882C820.806 309.305 820.236 309.899 819.797 310.664C819.357 311.429 819.032 312.316 818.82 313.325C818.625 314.334 818.527 315.425 818.527 316.597ZM858.405 324.385V312.202C858.405 311.307 858.251 310.534 857.941 309.883C857.632 309.232 857.16 308.727 856.525 308.369C855.891 308.011 855.085 307.832 854.108 307.832C853.246 307.832 852.489 307.979 851.838 308.271C851.203 308.564 850.715 308.979 850.373 309.517C850.031 310.037 849.86 310.64 849.86 311.323H843.391C843.391 310.233 843.651 309.199 844.172 308.223C844.693 307.23 845.433 306.351 846.394 305.586C847.37 304.805 848.534 304.194 849.885 303.755C851.252 303.315 852.782 303.096 854.475 303.096C856.477 303.096 858.259 303.438 859.821 304.121C861.4 304.788 862.637 305.798 863.532 307.148C864.444 308.499 864.899 310.2 864.899 312.251V323.774C864.899 325.093 864.981 326.224 865.144 327.168C865.323 328.096 865.583 328.901 865.925 329.585V330H859.357C859.048 329.333 858.812 328.486 858.649 327.461C858.487 326.419 858.405 325.394 858.405 324.385ZM859.309 313.911L859.357 317.744H855.28C854.271 317.744 853.384 317.85 852.619 318.062C851.854 318.257 851.228 318.55 850.739 318.94C850.251 319.315 849.885 319.771 849.641 320.308C849.396 320.828 849.274 321.423 849.274 322.09C849.274 322.741 849.421 323.327 849.714 323.848C850.023 324.368 850.463 324.784 851.032 325.093C851.618 325.386 852.302 325.532 853.083 325.532C854.222 325.532 855.215 325.304 856.062 324.849C856.908 324.377 857.567 323.807 858.039 323.14C858.511 322.472 858.763 321.838 858.796 321.235L860.651 324.019C860.424 324.686 860.082 325.394 859.626 326.143C859.17 326.891 858.584 327.591 857.868 328.242C857.152 328.893 856.289 329.43 855.28 329.854C854.271 330.277 853.099 330.488 851.765 330.488C850.056 330.488 848.526 330.146 847.175 329.463C845.824 328.779 844.758 327.843 843.977 326.655C843.195 325.467 842.805 324.116 842.805 322.603C842.805 321.203 843.065 319.966 843.586 318.892C844.107 317.817 844.88 316.914 845.905 316.182C846.931 315.433 848.2 314.871 849.714 314.497C851.244 314.106 852.993 313.911 854.963 313.911H859.309ZM889.055 324.385V292.5H895.549V330H889.689L889.055 324.385ZM872.087 317.109V316.597C872.087 314.578 872.315 312.747 872.771 311.104C873.243 309.443 873.926 308.019 874.821 306.831C875.716 305.643 876.799 304.723 878.068 304.072C879.354 303.421 880.811 303.096 882.438 303.096C884.017 303.096 885.393 303.413 886.564 304.048C887.753 304.683 888.762 305.586 889.592 306.758C890.438 307.93 891.114 309.321 891.618 310.933C892.123 312.528 892.489 314.285 892.717 316.206V317.598C892.489 319.469 892.123 321.187 891.618 322.749C891.114 324.312 890.438 325.679 889.592 326.851C888.762 328.006 887.753 328.901 886.564 329.536C885.376 330.171 883.985 330.488 882.39 330.488C880.778 330.488 879.33 330.155 878.044 329.487C876.774 328.82 875.692 327.884 874.797 326.68C873.918 325.475 873.243 324.059 872.771 322.432C872.315 320.804 872.087 319.03 872.087 317.109ZM878.557 316.597V317.109C878.557 318.249 878.654 319.315 878.85 320.308C879.045 321.3 879.362 322.179 879.802 322.944C880.241 323.693 880.803 324.279 881.486 324.702C882.186 325.125 883.033 325.337 884.025 325.337C885.295 325.337 886.337 325.06 887.15 324.507C887.98 323.937 888.623 323.164 889.079 322.188C889.535 321.195 889.828 320.08 889.958 318.843V315.01C889.893 314.033 889.722 313.13 889.445 312.3C889.185 311.47 888.811 310.754 888.322 310.151C887.85 309.549 887.264 309.077 886.564 308.735C885.865 308.394 885.035 308.223 884.074 308.223C883.081 308.223 882.235 308.442 881.535 308.882C880.835 309.305 880.266 309.899 879.826 310.664C879.387 311.429 879.061 312.316 878.85 313.325C878.654 314.334 878.557 315.425 878.557 316.597ZM925.28 308.662V340.156H918.811V303.584H924.792L925.28 308.662ZM942.248 316.523V317.036C942.248 318.957 942.02 320.739 941.564 322.383C941.125 324.01 940.474 325.435 939.611 326.655C938.749 327.86 937.674 328.804 936.389 329.487C935.119 330.155 933.654 330.488 931.994 330.488C930.367 330.488 928.951 330.179 927.746 329.561C926.542 328.926 925.524 328.031 924.694 326.875C923.864 325.719 923.197 324.377 922.692 322.847C922.204 321.3 921.838 319.616 921.594 317.793V316.157C921.838 314.22 922.204 312.463 922.692 310.884C923.197 309.289 923.864 307.913 924.694 306.758C925.524 305.586 926.534 304.683 927.722 304.048C928.926 303.413 930.334 303.096 931.945 303.096C933.622 303.096 935.095 303.413 936.364 304.048C937.65 304.683 938.732 305.594 939.611 306.782C940.49 307.97 941.149 309.386 941.589 311.03C942.028 312.674 942.248 314.505 942.248 316.523ZM935.778 317.036V316.523C935.778 315.352 935.673 314.269 935.461 313.276C935.249 312.267 934.924 311.388 934.484 310.64C934.045 309.875 933.475 309.281 932.775 308.857C932.076 308.434 931.229 308.223 930.236 308.223C929.243 308.223 928.389 308.385 927.673 308.711C926.957 309.036 926.371 309.5 925.915 310.103C925.459 310.705 925.101 311.421 924.841 312.251C924.597 313.065 924.434 313.968 924.353 314.961V319.014C924.499 320.218 924.784 321.3 925.207 322.261C925.63 323.221 926.249 323.986 927.062 324.556C927.893 325.125 928.967 325.41 930.285 325.41C931.278 325.41 932.124 325.19 932.824 324.751C933.524 324.312 934.094 323.709 934.533 322.944C934.973 322.163 935.29 321.268 935.485 320.259C935.681 319.25 935.778 318.175 935.778 317.036ZM948.312 317.061V316.548C948.312 314.611 948.589 312.829 949.143 311.201C949.696 309.557 950.502 308.133 951.56 306.929C952.618 305.724 953.911 304.788 955.441 304.121C956.971 303.438 958.713 303.096 960.666 303.096C962.652 303.096 964.41 303.438 965.939 304.121C967.486 304.788 968.788 305.724 969.846 306.929C970.904 308.133 971.709 309.557 972.263 311.201C972.816 312.829 973.093 314.611 973.093 316.548V317.061C973.093 318.981 972.816 320.763 972.263 322.407C971.709 324.035 970.904 325.459 969.846 326.68C968.788 327.884 967.494 328.82 965.964 329.487C964.434 330.155 962.684 330.488 960.715 330.488C958.762 330.488 957.012 330.155 955.466 329.487C953.92 328.82 952.618 327.884 951.56 326.68C950.502 325.459 949.696 324.035 949.143 322.407C948.589 320.763 948.312 318.981 948.312 317.061ZM954.758 316.548V317.061C954.758 318.216 954.872 319.299 955.1 320.308C955.327 321.317 955.677 322.204 956.149 322.969C956.621 323.734 957.232 324.336 957.98 324.775C958.745 325.199 959.657 325.41 960.715 325.41C961.757 325.41 962.652 325.199 963.4 324.775C964.149 324.336 964.759 323.734 965.231 322.969C965.72 322.204 966.078 321.317 966.306 320.308C966.534 319.299 966.647 318.216 966.647 317.061V316.548C966.647 315.409 966.534 314.342 966.306 313.35C966.078 312.34 965.72 311.453 965.231 310.688C964.759 309.907 964.141 309.297 963.376 308.857C962.627 308.402 961.724 308.174 960.666 308.174C959.624 308.174 958.729 308.402 957.98 308.857C957.232 309.297 956.621 309.907 956.149 310.688C955.677 311.453 955.327 312.34 955.1 313.35C954.872 314.342 954.758 315.409 954.758 316.548ZM986.726 308.979V330H980.28V303.584H986.384L986.726 308.979ZM994.758 303.413L994.66 309.419C994.302 309.354 993.895 309.305 993.439 309.272C993 309.24 992.585 309.224 992.194 309.224C991.201 309.224 990.331 309.362 989.582 309.639C988.833 309.899 988.207 310.282 987.702 310.786C987.214 311.291 986.84 311.909 986.579 312.642C986.319 313.358 986.172 314.172 986.14 315.083L984.748 314.912C984.748 313.236 984.919 311.681 985.261 310.249C985.603 308.817 986.099 307.563 986.75 306.489C987.401 305.415 988.215 304.585 989.191 303.999C990.184 303.397 991.324 303.096 992.609 303.096C992.967 303.096 993.35 303.128 993.757 303.193C994.18 303.242 994.514 303.315 994.758 303.413ZM1027.61 330.488C1025.61 330.488 1023.81 330.163 1022.22 329.512C1020.62 328.861 1019.26 327.957 1018.14 326.802C1017.03 325.63 1016.18 324.271 1015.58 322.725C1014.99 321.162 1014.7 319.486 1014.7 317.695V316.719C1014.7 314.684 1014.99 312.837 1015.58 311.177C1016.16 309.5 1016.99 308.06 1018.07 306.855C1019.14 305.651 1020.43 304.723 1021.93 304.072C1023.42 303.421 1025.08 303.096 1026.88 303.096C1028.75 303.096 1030.41 303.413 1031.84 304.048C1033.27 304.666 1034.47 305.545 1035.43 306.685C1036.39 307.824 1037.11 309.191 1037.6 310.786C1038.09 312.365 1038.33 314.115 1038.33 316.035V318.745H1017.63V314.302H1031.98V313.813C1031.95 312.788 1031.76 311.852 1031.4 311.006C1031.04 310.143 1030.49 309.46 1029.74 308.955C1028.99 308.434 1028.02 308.174 1026.83 308.174C1025.87 308.174 1025.03 308.385 1024.32 308.809C1023.62 309.215 1023.03 309.801 1022.56 310.566C1022.1 311.315 1021.76 312.21 1021.54 313.252C1021.31 314.294 1021.19 315.449 1021.19 316.719V317.695C1021.19 318.802 1021.34 319.827 1021.63 320.771C1021.94 321.715 1022.39 322.537 1022.98 323.237C1023.58 323.921 1024.29 324.458 1025.12 324.849C1025.97 325.223 1026.93 325.41 1028 325.41C1029.36 325.41 1030.58 325.15 1031.67 324.629C1032.77 324.092 1033.73 323.302 1034.55 322.261L1037.79 325.63C1037.24 326.444 1036.49 327.225 1035.55 327.974C1034.62 328.722 1033.5 329.333 1032.18 329.805C1030.86 330.26 1029.34 330.488 1027.61 330.488ZM1051.99 292.5V330H1045.52V292.5H1051.99ZM1089.7 314.155H1080.62L1080.57 309.419H1088.36C1089.7 309.419 1090.81 309.232 1091.71 308.857C1092.6 308.483 1093.28 307.938 1093.73 307.222C1094.2 306.506 1094.44 305.635 1094.44 304.609C1094.44 303.47 1094.22 302.542 1093.78 301.826C1093.36 301.11 1092.69 300.589 1091.78 300.264C1090.87 299.922 1089.71 299.751 1088.31 299.751H1082.79V330H1076.08V294.453H1088.31C1090.33 294.453 1092.13 294.648 1093.71 295.039C1095.3 295.413 1096.65 295.999 1097.76 296.797C1098.87 297.594 1099.71 298.595 1100.28 299.8C1100.86 301.004 1101.15 302.437 1101.15 304.097C1101.15 305.562 1100.81 306.912 1100.13 308.149C1099.46 309.37 1098.43 310.363 1097.03 311.128C1095.64 311.893 1093.89 312.332 1091.75 312.446L1089.7 314.155ZM1089.41 330H1078.64L1081.45 324.727H1089.41C1090.75 324.727 1091.84 324.507 1092.71 324.067C1093.59 323.628 1094.24 323.026 1094.66 322.261C1095.1 321.479 1095.32 320.584 1095.32 319.575C1095.32 318.468 1095.12 317.508 1094.73 316.694C1094.36 315.881 1093.76 315.254 1092.93 314.814C1092.11 314.375 1091.04 314.155 1089.7 314.155H1082.72L1082.77 309.419H1091.66L1093.2 311.25C1095.25 311.266 1096.91 311.673 1098.2 312.471C1099.5 313.268 1100.46 314.294 1101.08 315.547C1101.7 316.8 1102.01 318.151 1102.01 319.6C1102.01 321.878 1101.51 323.791 1100.52 325.337C1099.54 326.883 1098.11 328.047 1096.22 328.828C1094.35 329.609 1092.08 330 1089.41 330ZM1124.38 324.385V312.202C1124.38 311.307 1124.23 310.534 1123.92 309.883C1123.61 309.232 1123.14 308.727 1122.5 308.369C1121.87 308.011 1121.06 307.832 1120.08 307.832C1119.22 307.832 1118.47 307.979 1117.81 308.271C1117.18 308.564 1116.69 308.979 1116.35 309.517C1116.01 310.037 1115.84 310.64 1115.84 311.323H1109.37C1109.37 310.233 1109.63 309.199 1110.15 308.223C1110.67 307.23 1111.41 306.351 1112.37 305.586C1113.35 304.805 1114.51 304.194 1115.86 303.755C1117.23 303.315 1118.76 303.096 1120.45 303.096C1122.45 303.096 1124.24 303.438 1125.8 304.121C1127.38 304.788 1128.61 305.798 1129.51 307.148C1130.42 308.499 1130.88 310.2 1130.88 312.251V323.774C1130.88 325.093 1130.96 326.224 1131.12 327.168C1131.3 328.096 1131.56 328.901 1131.9 329.585V330H1125.33C1125.02 329.333 1124.79 328.486 1124.63 327.461C1124.46 326.419 1124.38 325.394 1124.38 324.385ZM1125.29 313.911L1125.33 317.744H1121.26C1120.25 317.744 1119.36 317.85 1118.6 318.062C1117.83 318.257 1117.2 318.55 1116.72 318.94C1116.23 319.315 1115.86 319.771 1115.62 320.308C1115.37 320.828 1115.25 321.423 1115.25 322.09C1115.25 322.741 1115.4 323.327 1115.69 323.848C1116 324.368 1116.44 324.784 1117.01 325.093C1117.59 325.386 1118.28 325.532 1119.06 325.532C1120.2 325.532 1121.19 325.304 1122.04 324.849C1122.88 324.377 1123.54 323.807 1124.02 323.14C1124.49 322.472 1124.74 321.838 1124.77 321.235L1126.63 324.019C1126.4 324.686 1126.06 325.394 1125.6 326.143C1125.15 326.891 1124.56 327.591 1123.84 328.242C1123.13 328.893 1122.27 329.43 1121.26 329.854C1120.25 330.277 1119.08 330.488 1117.74 330.488C1116.03 330.488 1114.5 330.146 1113.15 329.463C1111.8 328.779 1110.73 327.843 1109.95 326.655C1109.17 325.467 1108.78 324.116 1108.78 322.603C1108.78 321.203 1109.04 319.966 1109.56 318.892C1110.08 317.817 1110.86 316.914 1111.88 316.182C1112.91 315.433 1114.18 314.871 1115.69 314.497C1117.22 314.106 1118.97 313.911 1120.94 313.911H1125.29ZM1150.03 325.41C1150.94 325.41 1151.75 325.231 1152.47 324.873C1153.18 324.515 1153.75 324.01 1154.18 323.359C1154.62 322.708 1154.85 321.951 1154.88 321.089H1160.96C1160.93 322.879 1160.43 324.482 1159.45 325.898C1158.47 327.314 1157.17 328.438 1155.54 329.268C1153.93 330.081 1152.13 330.488 1150.12 330.488C1148.09 330.488 1146.32 330.146 1144.8 329.463C1143.29 328.779 1142.03 327.827 1141.02 326.606C1140.02 325.386 1139.28 323.97 1138.77 322.358C1138.28 320.747 1138.04 319.022 1138.04 317.183V316.401C1138.04 314.562 1138.28 312.837 1138.77 311.226C1139.28 309.614 1140.02 308.198 1141.02 306.978C1142.03 305.757 1143.29 304.805 1144.8 304.121C1146.32 303.438 1148.08 303.096 1150.1 303.096C1152.23 303.096 1154.1 303.511 1155.71 304.341C1157.34 305.171 1158.61 306.343 1159.52 307.856C1160.45 309.37 1160.93 311.152 1160.96 313.203H1154.88C1154.85 312.259 1154.64 311.413 1154.25 310.664C1153.86 309.915 1153.31 309.313 1152.59 308.857C1151.87 308.402 1151 308.174 1149.98 308.174C1148.89 308.174 1147.98 308.402 1147.24 308.857C1146.53 309.313 1145.97 309.94 1145.56 310.737C1145.17 311.519 1144.89 312.397 1144.73 313.374C1144.58 314.334 1144.51 315.343 1144.51 316.401V317.183C1144.51 318.257 1144.58 319.282 1144.73 320.259C1144.89 321.235 1145.17 322.114 1145.56 322.896C1145.97 323.66 1146.53 324.271 1147.24 324.727C1147.98 325.182 1148.9 325.41 1150.03 325.41ZM1174.21 292.476V330H1167.76V292.476H1174.21ZM1190.76 303.584L1179.26 316.499L1173.03 322.822L1170.98 317.817L1175.79 311.763L1182.97 303.584H1190.76ZM1184.17 330L1175.99 317.695L1180.29 313.521L1191.64 330H1184.17ZM1208.05 330.488C1206.05 330.488 1204.25 330.163 1202.66 329.512C1201.06 328.861 1199.7 327.957 1198.58 326.802C1197.47 325.63 1196.62 324.271 1196.02 322.725C1195.43 321.162 1195.14 319.486 1195.14 317.695V316.719C1195.14 314.684 1195.43 312.837 1196.02 311.177C1196.6 309.5 1197.43 308.06 1198.51 306.855C1199.58 305.651 1200.87 304.723 1202.37 304.072C1203.86 303.421 1205.51 303.096 1207.32 303.096C1209.19 303.096 1210.85 303.413 1212.28 304.048C1213.71 304.666 1214.91 305.545 1215.87 306.685C1216.83 307.824 1217.55 309.191 1218.04 310.786C1218.53 312.365 1218.77 314.115 1218.77 316.035V318.745H1198.07V314.302H1212.42V313.813C1212.39 312.788 1212.2 311.852 1211.84 311.006C1211.48 310.143 1210.93 309.46 1210.18 308.955C1209.43 308.434 1208.46 308.174 1207.27 308.174C1206.31 308.174 1205.47 308.385 1204.76 308.809C1204.06 309.215 1203.47 309.801 1203 310.566C1202.54 311.315 1202.2 312.21 1201.97 313.252C1201.75 314.294 1201.63 315.449 1201.63 316.719V317.695C1201.63 318.802 1201.78 319.827 1202.07 320.771C1202.38 321.715 1202.83 322.537 1203.42 323.237C1204.02 323.921 1204.73 324.458 1205.56 324.849C1206.41 325.223 1207.37 325.41 1208.44 325.41C1209.8 325.41 1211.02 325.15 1212.11 324.629C1213.21 324.092 1214.17 323.302 1214.99 322.261L1218.23 325.63C1217.68 326.444 1216.93 327.225 1215.99 327.974C1215.06 328.722 1213.94 329.333 1212.62 329.805C1211.3 330.26 1209.78 330.488 1208.05 330.488ZM1231.92 309.224V330H1225.47V303.584H1231.53L1231.92 309.224ZM1230.89 315.84H1228.99C1229 313.919 1229.26 312.178 1229.77 310.615C1230.27 309.053 1230.98 307.71 1231.89 306.587C1232.82 305.464 1233.92 304.601 1235.19 303.999C1236.46 303.397 1237.87 303.096 1239.44 303.096C1240.71 303.096 1241.85 303.275 1242.88 303.633C1243.9 303.991 1244.78 304.561 1245.51 305.342C1246.26 306.123 1246.83 307.148 1247.22 308.418C1247.63 309.671 1247.83 311.217 1247.83 313.057V330H1241.34V313.008C1241.34 311.803 1241.16 310.851 1240.8 310.151C1240.46 309.451 1239.96 308.955 1239.29 308.662C1238.64 308.369 1237.83 308.223 1236.87 308.223C1235.88 308.223 1235.01 308.426 1234.26 308.833C1233.53 309.224 1232.91 309.769 1232.4 310.469C1231.92 311.169 1231.54 311.974 1231.28 312.886C1231.02 313.797 1230.89 314.782 1230.89 315.84ZM1271.87 324.385V292.5H1278.36V330H1272.5L1271.87 324.385ZM1254.9 317.109V316.597C1254.9 314.578 1255.13 312.747 1255.58 311.104C1256.06 309.443 1256.74 308.019 1257.63 306.831C1258.53 305.643 1259.61 304.723 1260.88 304.072C1262.17 303.421 1263.62 303.096 1265.25 303.096C1266.83 303.096 1268.21 303.413 1269.38 304.048C1270.57 304.683 1271.57 305.586 1272.4 306.758C1273.25 307.93 1273.93 309.321 1274.43 310.933C1274.94 312.528 1275.3 314.285 1275.53 316.206V317.598C1275.3 319.469 1274.94 321.187 1274.43 322.749C1273.93 324.312 1273.25 325.679 1272.4 326.851C1271.57 328.006 1270.57 328.901 1269.38 329.536C1268.19 330.171 1266.8 330.488 1265.2 330.488C1263.59 330.488 1262.14 330.155 1260.86 329.487C1259.59 328.82 1258.5 327.884 1257.61 326.68C1256.73 325.475 1256.06 324.059 1255.58 322.432C1255.13 320.804 1254.9 319.03 1254.9 317.109ZM1261.37 316.597V317.109C1261.37 318.249 1261.47 319.315 1261.66 320.308C1261.86 321.3 1262.17 322.179 1262.61 322.944C1263.05 323.693 1263.62 324.279 1264.3 324.702C1265 325.125 1265.85 325.337 1266.84 325.337C1268.11 325.337 1269.15 325.06 1269.96 324.507C1270.79 323.937 1271.44 323.164 1271.89 322.188C1272.35 321.195 1272.64 320.08 1272.77 318.843V315.01C1272.71 314.033 1272.53 313.13 1272.26 312.3C1272 311.47 1271.62 310.754 1271.13 310.151C1270.66 309.549 1270.08 309.077 1269.38 308.735C1268.68 308.394 1267.85 308.223 1266.89 308.223C1265.89 308.223 1265.05 308.442 1264.35 308.882C1263.65 309.305 1263.08 309.899 1262.64 310.664C1262.2 311.429 1261.87 312.316 1261.66 313.325C1261.47 314.334 1261.37 315.425 1261.37 316.597ZM1286.96 326.851C1286.96 325.874 1287.3 325.052 1287.97 324.385C1288.63 323.717 1289.54 323.384 1290.68 323.384C1291.82 323.384 1292.72 323.717 1293.39 324.385C1294.05 325.052 1294.39 325.874 1294.39 326.851C1294.39 327.811 1294.05 328.625 1293.39 329.292C1292.72 329.943 1291.82 330.269 1290.68 330.269C1289.54 330.269 1288.63 329.943 1287.97 329.292C1287.3 328.625 1286.96 327.811 1286.96 326.851Z" fill="#3BA9C3"/>
<rect x="-0.5" y="-0.5" width="1377" height="477" stroke="url(#paint1_radial_367_2)"/>
</g>
</g>
<defs>
<filter id="filter0_b_367_2" x="-43" y="-43" width="1462" height="562" filterUnits="userSpaceOnUse" color-interpolation-filters="sRGB">
<feFlood flood-opacity="0" result="BackgroundImageFix"/>
<feGaussianBlur in="BackgroundImage" stdDeviation="21"/>
<feComposite in2="SourceAlpha" operator="in" result="effect1_backgroundBlur_367_2"/>
<feBlend mode="normal" in="SourceGraphic" in2="effect1_backgroundBlur_367_2" result="shape"/>
</filter>
<pattern id="pattern0" patternContentUnits="objectBoundingBox" width="1" height="1">
<use xlink:href="#image0_367_2" transform="scale(0.00239808)"/>
</pattern>
<linearGradient id="paint0_linear_367_2" x1="0" y1="0" x2="1090.99" y2="844.291" gradientUnits="userSpaceOnUse">
<stop stop-color="#158AF6" stop-opacity="0.3"/>
<stop offset="0.385599" stop-color="#5062D8" stop-opacity="0"/>
<stop offset="0.483825" stop-color="#595BD3" stop-opacity="0"/>
<stop offset="0.599613" stop-color="#6553CD" stop-opacity="0"/>
<stop offset="1" stop-color="#BA1AA0" stop-opacity="0.25"/>
</linearGradient>
<radialGradient id="paint1_radial_367_2" cx="0" cy="0" r="1" gradientUnits="userSpaceOnUse" gradientTransform="translate(688 238) rotate(161.194) scale(738.299 1076.67)">
<stop stop-color="#151515"/>
<stop offset="1" stop-color="#151515" stop-opacity="0"/>
</radialGradient>
<clipPath id="clip0_367_2">
<rect width="1376" height="476" rx="20" fill="white"/>
</clipPath>
<image id="image0_367_2" width="417" height="417" xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAAaEAAAGhCAYAAADIqAvCAAAACXBIWXMAAAsTAAALEwEAmpwYAAAAIGNIUk0AAHolAACAgwAA+f8AAIDpAAB1MAAA6mAAADqYAAAXb5JfxUYAAbo+SURBVHja7P13gCzXdR6If+fce6uqw8SXAx5yJggCDKJIihQjGMUoUiJFWmnX2uCw3rV3LXvltaxoSrLlIHnt33ptWZYtr0SJli1ZokRSjCJFEAQTQBI5Pjy8NDMdquqG8/vj3uow0/PeA5NAog7YnDcz3dXVPdX3u+ec73wfiQjaaKONNtpo4y8iuH0L2mijjTbaaEGojTbaaKONFoTaaKONNtpoowWhNtpoo402WhBqo4022mijjRaE2mijjTbaaEGojTbaaKONNloQaqONNtpoowWhNtpoo4022mhBqI022mijjRaE2mijjTbaaKMFoTbaaKONNloQaqONNtpoo40WhNpoo4022mhBqI022mijjTZaEGqjjTbaaKMFoTbaaKONNloQaqONNtpoo40WhNpoo4022mhBqI022mijjTZaEGqjjTbaaOPbN/S34kkTUfuX2yWefsWNuYgUAskAmPg3FgURBSKBACB4AB4gRyBLRJZA5e13faZq38Enb4hI+ya08W0X9K14YbcgBDzj8hs63rt+EOkz8zKAZRfcmg/+AAgHSfEeIloBU5+JCiEyLCAhCSSovcgIIQwA2hDrT4Ho0cLkx5XSZ0joNIANYrX5qS/dWrYfkxaE2mijBaGnOAjdcNnTtEhY8+L3QMJBH/ylLvibSOsrTZ6tK6X7YO6wUhkrLpjYgEiBSAFQICIGIf0viMAD4kXEIYTaeV/B+zGATQrhRF3Wd3LAn2tl7mKix4no1Ke/cvug/ci0INRGGy0IPUVA6OmXXdez1q5Ya/fZ4C/WhX6+ysyNpNUhIdpDUP0szztam2zR31HiygViBhOBJjcG0fR9JCKEECaLXAjB2roautqeEe+Pq+C/BCvvh9Anmfixz973hbPtR6cFoTbaaEHo2zBuvOz63Dm7x9r6IkG42iG8zBNfC6P35kW+orOib4wyBAZAYFYAZLJAicjc+0Nz4ENg5jnwAQBmRghhbqFrQCmEgGo02ArOPe7L+k7Y8F8Z/BGt9QOff+DOFoxaEGqjjRaEvj3A52lLVVUedK6+RhRe7UmexcYc0nm+pnTWZaXArEFE0EZDsYL3DiGECcCITMFoFmiYeSEgNaGU2rHQzYIQQoBzFlVVVbYsH7fj8svKy29nOvsTo83Dn73/jrZM14JQG220IPStFjdfe3PurN3nnT1W1eX1tbev10Vxbdbp7DXGLMcyGgPEIB2Bp8lcIkB4iHgA8wC0HYSUUnPfLwKiWSBrFrwGhDQzrLWw1sJ7B+dcXY1Gx0NZ3mrAv6V19gmt1cOfvffOlsTQglAbbbQg9GSPm669qe+cOyTwN1pvX1IH/x1Ft3+Ild5rjDFKKxBxAhw1ARkiTsAjE8BgJsyW47YDzaL3bfvvZ/89W84LISCEAO9DLONJgHMO1lo4Z1FX1cjX9aPk7J/pwP9Gm+xzn7//S4+1H6sWhNpoowWhJyP4XHdz3zt3zPv65lrcm8mYp+s835eZfIlZTQBg2rehyVcRAhEgEibZUFMyY46/222xmu0DLXoPZwEoHi/e33sP7z2YdQQ67+C9nwBUyopg63LTleN7tcdvZip7r9Lm7tvv+WI7c9SCUBtttCD0ZIhnXv9ssrY6WrvqmaT5HZSZZyqdHTTGdJjVhLE2XWho24JDABhEAkDmMhgRgCg8ofdrUUY0+3wNGE1Lcw1IBYjE7EiCAJPvPeq6gq3Kh9n69+ug/pU22Wc+e+8Xt9qPWAtCbbTRgtBfYNx87c0ro9HwUgf3LmT6Nb2lpSNK6x7F0Z0JaaBZ6BcvNruDUHpEuj1xENr+++09oebcpv+OoCMhAJPzlGmZzpZnw7i6VXv6p8bkH//8A1860X7MWhBqo40WhL7J8ezrbs6td8cCyYsH1fitvaWVG/JOZz8rBmS+9xIX/O2vibe95u2kA5qA0hN9385VmpsFoe3nFv8dIOIRQgIpEVACRudcKhGGshoM77aD4a93su7v5EV+7+33fLFuP24tCLXRRgtC34R45tU37q1teZMo/JDu959riuIwQeUNq207ky3+m7ctMrytbxMWAMk8HXu3v2UDeE/kfZs9VhohmgGhMMeeQwgwxkAkwHs/6SeNh4Pjfjj6UKHyX8mL/LOfufuLZ9qPXAtCbbTRgtA3Kvu59ma2tr7YhepV1O38oM6Lq5Uxy0opSFi8mMyWurZnQlOgkQhCRKCJ9M6Fvwezs0RPdMGbL8vJjhsAqJm+UsOoa8LZaqsejr6ovfyLTlb88W33fPGh9mPXglAbbbQg9HWOm6+6ccXW1fWe3V8yvd4riuXli5iVahZmmimvbS91bVc5aEBo+lo9gBDBZzYTErqgBWvR/NBu7+ficpzs+j0AaOYJa26W3t3MMnnvra/Ke7ULv5Gx/g/a6Ls/9eXP+/bj14JQG220IPR1iBsvf/oB68Yv9kr+u3x5+RlZ0Vln5gnpIIQAJrVrhtGAzuJynCQAims2s1qwOu1OalgERufqCZ0PeLaDVERGhngPFgIrnmZF4uG9m5TvXF09yJV9b876X2mt77j1ri/Y9iPYglAbLQi1IPQ1xHXHrr3Ehfq1VOi/rLvdK4tOJzfGAEIQBEBoR89mdkGfUqR3IyY0IDSdD9oNhHbLfrY/9/nYcU8kC4rMPQITgQXwYdq7CuLBHAGprit47xFs/RjX9g9zNr+cZeYLt97VzhO1INRGC0ItCD3huP6Sp2lbV1cH8t+HIntH0e9fYowhrTVYq5TZ+OSkEEACgGYW8B29oJ2Z0BwILaRm775QzYMFP6H3c2fvx+8AuFnV7e3qC4vOSUTi8KuzsOX4FKr6j3qm+OXcmNtvvfuLrdxPC0JttCDUgtCFZz/Xdcbj4Q1O3A+rpe5ru/2lI3negVIKrNXM7E+zSAsQBJihWZ8PhJrMqCnJRY04Oedsz+6ZD2O3P/O5QGMWhBb/XHYFoNneUBPee4iPJbpqPDpFtf3jvil+MTP69k/fc2dL4W5BqI2nYOj2LXhicc1F13RHo60bLbn/1fS6Lyw63X1aayilolAo84JFPmm9bZvp2a5UMP99QFROQAIhbAOTWfBYRDZoAGj6/TwwXhiQN6oMu53z+UBtuy5dvDF0lu9xwEtKVw0J8ksAvtBeXW208dQLbt+CC49rj12bjUeDp9dS/01V5C82eb5PKQWtdRISxa4NfEFYmG3slr0sOta5sxVZCAjnEis93/0X3XYDsN08jBoduok0EcV3AwBYm32W6ZbSVd93/ZFLL2qvsDbaaEGojV3iuouvo7oaX+HJ/6jq5N+lTLaulYI2BlrrifYbgsxV3WaVDiJ6LKZWx5LXdg24ph8TFgLPE41zZT/nMsKLl8n8beocvvhnzb+Z1QyZogHXaQYnSh+pWN5ivXvB045ettJeaW200YJQGwvC1tVR6+s3cWFeYfJ8r0oApJRKfY/dmWlPFEAW9VYuJL6ePYNFmc+FZEq0w0Z8/rUwReo6M0OpNAtlsksruB+t6uqGp110mWqvtjbaeOpE2xO6gLjm6FVrVTW8Bbl6p87zi5goMuDSIhqlatScnQKlhnyYaIzKbDJwjggTGZ9ZYLmQPsy5ymznA6jtA7Pb77+of9X87Fxlu6an1BAUiKclumgboSAiedD6GVVt30bWPQDggfaqa6ONFoTaAHDt0at0VY6e5lT4YTb5ZSIC0k0fKPY4tEp+O7Pkt6aENvl5I8B2fsWCWNoLEGnAINo7nOtxX0ucS3PufKC2HXRm55ji74DGF4mIZ2txEzmhEAJI6XXR4RZb1R+99tDFZ+949P7N9upro41v/2jLcecJa+t9jvzrOc+vJiItxCBlwCopICSttMZqe3pLOmo+QEKAd+mWjOK89xOdtanEzfRYITQ9ohkPn/MoGSwChtmZngshPCx67Ln7RfOAOD2HxSzBRdlUk02KUse8wrtq566+7sil7bXZRhttJvTUjqsPX5kNBxs3Ske9yii1LiKg2UU8ZTnb1QguZLE/V+ax/ThTh9XZRX1xFtVkTdMsZBHbbvKIuePPUrpnf9+U0mY9hRad1zxAzWZMO1mA21+rUhoh+LwG3YzgXsdOPQqgFTtto40WhJ664azdB0Vv1ln3IgmCQDJNHYWAQBCazxZmlQQulD59YSrX88cIoZHwmT9OfCpK4BjSfBFt6y017q3x90pN548aUJ0MowIIC9QSAMxp4zWluKbfM6+dl/pGzAjep+fARFNuysATsMkOeHKvC8Anrj1y6ck7Hr63VVNoo40WhJ56ceXhK/NyOLgBhX4Ba7XkvAWI4jwQYded/ez3IYSULckOQsJuTfx5t9QIKM3vzzdXtFOjLv2bYm8q+ICQFn4kEAgiYM+QILuW92JpcGrx3QBtM5wbbSViL2vKfIvDu9vPN4SQQE1iOpeGaufyJa0vLav6zQTcAeCe9mpso40WhJ5yEZxdJ8OvJZMdni7CKfMAnbPMNtvfkcR2k7A7CC0a7hTMSP6AtpEeZIcKQSqOzQHk/DkEeB97UgKBhGmvqAG4xSrZCSuI544JAEHCTAYmMxkRgTmCkGIFTRyVJETgQoAPIdI0iAAGgg/wkgA7nv9KYLwggzz72iOXPXrHw/eM2yuyjTZaEHpqleJcfQky9TxWajlImFmMabIAs/BCV9PZBb3JPIKXhQDUuK1GxYVURovpwVx2s71XIwB88FPgEUEQSbbbASHIhPzgvJ2Ax/ay37kYcNuBdbbMNkvNbr6f7R1NBUs9Kh9mwLWx6WvM+mhqEz4DhlDqSOnqNyivPgXg7vaKbKONFoSeQqW4K5ZsPX6WJxykCQlhmmRIWvB3k97Z7bZb1iQCNGQygczRmKeZyjZwmCFHNJmZ8w7eReDx3u9gxm0HkkWgs5ui9jwNm7CIMq6UWviamWZszZuyW1IUb+SOtgObEHUrWz+nA3nOdUcvf+iLD93dWj600UYLQk+NsM6tWPHfGVivcUpDpOlhJKCgGRBIPwQmbLkwc9sNhKKrKmheJPRChkpnS34iAufmKd9Ii31iJcypes+CyfZS3KKBVABRlggUB01T3yf2giZCPNP7C1JG5hFCAtSASUYos+BGiTiBKabNgiArfagO9rXK4eMA7muvzDbaaEHoKRHe+xVRdBlrVUwb5jMkAiT6M8mErjxZwCeNdpn2gxYYykXCQgQMzXqGBBB2ZcnNzxKFCfB4P589RXmcGYDD7mW4JgNpHrd98JSIoFinnzGYaeYrLTzubPbVnGPz2uZ/z9sypzA5HxGBybKOr+tnO++fe+3hy47f8cg9LVOujTZaEHoKBMkeKLU26WFcwJjPoob+LN15yi5rFvxJQrSjVLYoG9k+5DpX7lIMhtpBWJiCA8/1s2YBZzs7b5ZiPflZsibf/vPtwLWojDf77ylo+gUDusm6An4CjgAgSh2y3r/G+HArgK+0F2cbbbQg9G0dlx++IvehvigoWmLmuWb+dn213UBoYfmNZkjIJHN23rPZz6LHNwv4bPN/ulA37Ln552sW8TifM9/L2aF6QFNmHRPvBCjwDuDarYe0vdw3+xqa91NrvSNbmtwCz9HAA6s+ZfTC2ro3XXfkin/zxYfveqy9SttoowWhb9sI3nWI5Vpi1ZvPXOjrqNU2bzLXzNzMLsq706VnshlQ04raleo9yZQmGUwDOOm+2DaRlH42+wuBXJAI6rlebzNEu1PcdJ4swSEOtHqKckfgAGXMYaH6B7z4jadddOVvf/7BrzzeXqlttNGC0LdlSHAdMC4nRmeRkvR2kc7tILHo/s19pgSE7cOl8zbY28tti48dLcCJFFhtK5+lYdFFgLQoa5koXG/Pbp4A5i4C6e2OrJE+vtjQb/Y8AzHgPAI8WAtApJ1WV9Qh/Jh4p68/csXvsFaPfO7+L7V+12200YLQt1kmFHxfQIdEYETC3EI+u5hvH/DczjZbAG8LLLYxASXv50Ftke33dKFPQMM8MY3bngXN9252nvNsMKvFIDQ5n7BQrPR8fSGaKTtOdema81dzZn3b+2FaAyEQRCVZI88FjL7Gkv0rthpdnIX8d6+/6Mq7lFanPnvvna69cttoowWhb5dUaB3Q65BYhtpuTXB+ENvpgtosyNMa12wBTBCVss9tud3I4CilUt+Gd4DPbgrX82LpaVR0F0bc9tc5O8sz+7Pt99kuHbQInKYEDQUiP8mWtltDzJIjfACUMeDY98qF6CoL+cEq+O9yzn20QP4HT7v4qs8TqxOfu/eO0F7AbbTRgtC3dDDT3lrCMp+31CQLF+HdrAq2g8yUqryYfTervxZvekK9ns1uZp9neo6USnWYK/8toorvltlse092ANBux9ou99O8vvkMsVHyjr5J5wJfQcz0VJ5HuZ/gQVrvFe/2eGuvHAf3oizwHyqR33vaxVfd/fn7v9z2i9poowWhb8248tClhQ/VMRC6mFnwFykMzGY958qSmsV39r7zTLqmPDVVDmBmaK2hVDTPi2ZwsxQCLATE7V4+ISwWNl30+HOd//nsYHc7bnx+Tq9Rtomz8szzzlPY5wZWKQqkRg8nQZBEUweIiNedc2uVhKNiq+9SQf7rNYcv+y9Kqfu+8OBXhu0V3UYbLQh9S4XzPg/ij7A2WUw2FtORd+v97OYlNA9CDU16mvE0oZSCVgZaK2htkhAoJz25nbNGO4GAdpAfzgUcizKYRRnS7LHOpea98zliGXLnMXnmmI0dhexKWJh+jYoMBELAhD5PIYQDnniPtdVldT16Vu7Nr11z+NJP3vnIvS2du402WhD61gnvvQkI+wNgeKIns3sPZJGb6W4gNH34YvtrpRhKaRhtJtbh55LUWQQczUJ9rtLhPIhOfvJ1oZ+fj5CxKGvcbrC3SDpoLjMCQxrVBhEoZjhnAYgmyo84UreMqtHlurb/6coDx35PaXPXnQ+3unNttNGC0LdABO+Np7DGQnoGgxYutLuJl+4OVLwjm0rwA1aMIs/B3GRAjHkSQzhPZkNzXxfp1C06v+lCzzOkgcVAtuMZt5EJduuJbRdAXQRE8XG7ubtuf16e/D4ESeXLeM7eWwC0RNy9UZzdZ717Nlz4jasPXfKxLz1636PtFd5GGy0IPblBSMQIowsilQwVdsz6bAeZ7Yvq9hLc9kxpMkCaFk8mDa01jMlS/0nNEQym4BO2ZTHby1x8rhxl29ftwBp2ld5ZBBi7gdGix28Hq92BiHe8zkWgPbs1YCaI92BWyDKC9wxrLQCwMB2VIGvW+6vDuPytK/Yf+02TmXvuaNW422ijBaEna4iIBigHhM9Xatq+w1+kbj27SM+pAjCDwFCqISDoNKtDCzKbMNdHWbygnztzmSUGXKjqwfnICotKhLv1qiLNG7sC0fz80k5171mQ2v4cLkQrC0UEKD2jLO4gQA9KXU8ds+6su5Is/vm1Ry///B0P3b3ZXu1ttNGC0JMShARi4kq4+45+Udlpu2/P7ALbsN0aMdCJOrVS0FqBWW8bGCUs0oPb3h9pmGVECouKh/MLeDjPMO1CuNkV+M5FzNiRxVD0X6IIvZM+2PbSW2ODMQfqybBvmtPJ9NsgUMogBA8bHBiYsRSPFhcSHAKrQ8jo1fBhH4n/lWuPXv6hOx66+3R7xbfRRgtCTy4QCkI+CLMIFAAK0Y6BCSDWc144TflL0n0E83bZDchM7RAUiBlMOlK/0xwQJ9WDneWz2QWa5qwX5hf+pp8ju5ThGOCUSSUDPVBYWK1r6OJTll2a4+HGC1XmC2I0c65A9FiaWnTHxxAlxz6CEBDAoDQ3FMluMnFWnVK1JYq8AgiNknmYiiKE9HyAgCTp7FEcbIWE+KpZQymCYyBYB1J61TGeF5xdyoLk1xy97H13PnRPC0RttPEXHNy+Bdt24kEWCKDRDifVeeIBdpTgmhkfrTW0MmA2YIqzP9woHyQCwoVkJosqY9tlcxbbM8z2Uui8KuDNZSFCO17jJEMDxRRl9gaCEEfQmSE4TMz1IqJMHWEbS+90r8ZPCPMpKBBCvEmAFw8JHiQBEnxS2/YICYhC2gwgKYFDcQTAhujB3JMsu9Eq/HXr3UuvPXrpWnvVt9FGmwk9GctyOwEHfgcSNJv3iUV3IhbMAtAUGNSuGnTbS36Ly150TqrzOXcajX4bABE/sQNHA1A0k2MITe4PAIEEBI50AZlSJXgGHZtsJh5NpQwoHp5FALhoshfHTuMTBkpDuPF5SfwEjNBYnIuAwwxAEcABCAjpvpiW7BDikRnJWVbAArBEjT2JaRIUo0OZeXqQ+q/74Nz1Ry99/xceunejverbaKMFoScD/AAisgiEgsTSEm9jwUHmlauVUjDGzJXioqGcnstUdpO9WZwFNb2Z+Z+d73E7ezZyzsyrAYAgM+AIQHxMYliAwASW+eLfJEtqXlMU3osWEBAwBEi9nsj5aHpeIVUJp3p2k3No1B6a5EgmUDgZbCUECG0X/0lgzQIlDASAmOFDshwXwBjdRZbd6Ovqr3Jwo6cdvfSjn3/o3kF7/bfRRgtCf9EY5EXEL86EUk+E1Lbme1ywsyybk9qZSv1QYoepOQvveVVsnDMbmltcv4pQNPNaJtnL7vNEoDCVWA0MYZkkTfCyo/s0OefmNcwBVECQMKMgnhxUm0zQR0WIMKnaUezrpHIgT5OiSG6gKXkhyNSeXGgbzZwVEARaqZi1+SbDAoIVMKNHWfZMV1d/jbzbvP7opbd94aF7W/vwNtr4JkfbE5pfTb2I2BCCzFKtp1kPdgCQ4pj5NLcsM5NSXEM6UErvqqSwW/ay/X7nesz5MqDZ0t18v4jPqQQxKUN6F4kB6SsFH8t6wac0afqVEEASAPGgEJKBHqd8iKd9I4k5UhCBlwAfQhIoDfABsMHDeY86fXXewwek+wE+NGBOEw2+6U1BAk0ub1YKitWcBmCscKolMea5juV/Ct5ffv3Ry9vPQxtttJnQXyAiE3kIagA+zgzNLPzUWC6k0hOiD48x2QSA4iKnZxa6KWtNxM+X8TA9znZ69SKcWZQx7fb99jke36gRYNoDEvETrtv2UdZZEIuvxEdGW2P0LVNiXNPpmZM4SiQ3SmUyL4sp5JPWT4glwPh2TXtAXgIgDB8LdOm5wyQrEwDBB8z6JTGbKXMRPrEbI0mBoACR9Jj06sisOSUvRXDHlff/DMB97SehjTZaEPoLAiH2JBhLCB4qvjfTjGCa/cwu9lpr5Hk+0/+ZAtB2t9TzWSY8ocqhXJjeW6MRt3NGiFNpy5/z8WECRJGI3giIzhXwZNokmsBqiOQEHwg2xDIahbCN5i2JuBBAEvtHCM1758EICGAwRRo8RKCmfPLUX/KRBEEMEhVJF6nMGShuHgIlqncqQ0aKd+rvCQFsDjqFN4pzj1x7+LJfv+ORe060n4Y22mhB6JsPQkyehIYAfAMcSqk0vjIvqaO1RqfTQZF35iy/d/aTmnxgdykaEZkZsjx/iW2RLffuZbpmTqfpB6Vjpa9xkDTMaMdhypprmGnbpHdCIg6oifrDvFJEk8lICBBSgHDs3yQSgQSPENx01gcBLPGYFGIpj8UjxGIgiGlHiigikBDLb0oZhKbvZRQIHt4DwgFkOFK4GRG0ErXPSwB5QCsNpQQOOBZA7xQfHrn28GW/f8cj97SqCm200YLQNxuE2JLDwHnnKMnoEBFYz7uYaq2RZbEM1xATpovvdjHPWduCnVlMc1/v/Xkzmu2Acz6foG2vbm4OZ1ZYValUtvMRHBDmAc8n9FLM4AbEROC8T9lNokfPKWJHR9YQPNjZiToCJ9BRiIQJby0QHIAAJoFqrMtVnO/xDasuTIE9QOCdRx0CQAoheAgUghB88GCtoVUs49nawuRxRivAIwRBSJTtIAnkBGDFOgR1eeWqt2vvv3Tt4cs+d8cj97S24W200YLQNy8Us1NKnXUirslOJs3stPhrpZFnBYqi2Nb7mc4LzYOQny1czQHJbo6k5y6tya7H2O04IgGeQhQ+mL1fuq+t6nScAE4svBDieXsReCgADBcCFM0M5HJi7IWGQp6GRiVMejdaAkwaMCWKj1eJ0KEpoLtSoDBddPIM3U6OTl4gz6YzVrlOfZwJo1DBBo+yshjWFltbA5za2sKZzRHGtYcVC40M1gHOeagih9gIYM7H98sYBSKdBlxjKVGzhjK0FJW37Q+Qdf8UbX+ojTZaEPpmBjE7xeqkiK3jYmUmIBREwIqhZ0gIjWbc+cpni363HVAupL+zCIDObzAXF1oSRBkeCpAQbeEaCnSmdCx8hZi5RIDyk4WfGRCK5IQgMukRNTM+3rs4C4QAhkA32QwTCgYKYmRGI88z9LoFOnmGIjMwmmGYYTSjkxkUWYYiy6AbHT3xUMSQxJprBmK9BJS1w9halD2DfWtdDEqH0xsDPH5mA5WrYZhT/yjEGSEQFIVEb4jZXwiA95HBJ1AACdiYg8GH14mX+64+cOw3vvTYA6faT0YbbbQg9M0BIeIKQo9BpJ4td4UQEABkrJFnkYQQQlgIRBeqDbq9JHe+TOiJgNS5AAkS4oBtavQ3skTe1/DWQcTHZZoTIYEA60ooZqgkA0RJf45DUiVggU6ZkVEKRmlkmUFmNHqZQi9X6OQG/U43glAnZjtKxUxHgcAiUaNvlukGQHyIBIVtdPk6d7AhR+Ud9gWBFcbGcIzjj3dxenMLZwZDbIwq+MCoA0EZg6AVaudhfQ2wShT1xGAkP3kvyGTHnFRv0yF85trDl3zijkfuq9tPRxtttCD0DY+7H7/PHVk6cEYrVc9K7oiE6HqaZVBKTTKQBojmS3IX/nzyRO68S0Z0IceURIzgxISb6o42tHOBhkAxJdkeAGgyoYAOp76Jj0OhOmU2mWZoImjFyI1GL8/R63aw1Oui3++hW3TQ72boFAqGk3W5IjAHUEDKujxIJJYBMdtXilH71C9iQLyPg68AcgUYBfQ6HYysgw+EXm6w2u9hczjA46fP4sTpAc4MSjy+sYm6qqCKPBJAFMOLwImPpAeJBnnUqHoT5UHxdS7UP0wexwF85cmxSaL2Q/otFr/4g28wvSJbyZj6GtQJIYgXGtgQTv/Yv/r/Rl+X5/iBN/D/+uu/G76Rr+OrXasu6Lr+Rh78W/HDeGz18EtdLr+i8uIqIp5M5Od5B6YoYLRZqPvW9EMu5Dy/mvf8XAOo5zweyTz4YGaWR2LJy1kLQKBShiPBgzhmahkBHQUYrZAbg16RY3V5Gatry1ju9dDLc3S7OQwTDBM0MTQzjI42FY2EDzPFXlFCGQmC4F2UQyWagFDUK40lvhACHCRmKyKAd1H0NAiQyoaVdWBlAKXhBLAuwIrAB8KwCrjn0cfwwCPHcWZzhFoCalaANrBCqH0AWEc1Bu8jCIYIdgAgrn5AO/erRpl/feejD7S07TaeGDi863v6h/au3nzpRUd/rJvnh8vR2Jg8Z6X06PhjJz9x30MP/XsruPN//te/7Z/osf/xu960v9/JL+0W5spOp7h8NKruPTMsP11b3Ps3fu03hy0IfYuC0JX7LlfDcvhmvZL9AmlzUQiSMh+g21mCMhlAmMmGYqbQiHUuOsfJ1xDmPFK322Ev/DtI+j+aszfCvJ3djK1BmP1lslgQAYuFSuZ480Omka1mtIZiQLOC0oRca/T7fSyv9LHc7WClmyFXKkoTKYYxGkWmoUmBmZArglKpXCchioUmqR4RQqD4Bk3JBQCDU4aWSpEhRGAKmGjyBYpqCpHl7iEhJJUGAXyA934iDmu9h/dRQduFyNzzojGwHo+eOoWTZzdwYnMLpwdjVIFQM6P2DCiDIJHEkNpcCRwJhOBh69szL39HKfOBOx65r3VlbeOC4ufe9upi72rxnKOH9v24Z/Msomy91+lS7SzA2gZfPz7a2vjUeFT+6tmtwUf+x//nPRekXfizb32V3rO6fNPBg+s/QqyuJZMfCpCuFxkplT04Pjv+08cfe+w9o9H4zr/1n/7z143d+Y3EibYcNxNBZE0Yzw7gpYZJRiTIUh9IUTPgmWZrKDSC0Nv0j5rOBoMbgVPFcC5eE4oJLu30hSllW43Ap0CSfMBUWIHhk7lbzBqSgGciCSiWKJUTfOrd8KTnoxkolMCwj1mK1uiYOOPU7XaRZwZL/T6M0ci1htbxPplRyPMceaZRaANNDFY8oaQj9WyitmqYGVZlQEX7BYk1wKbLA+aZzBGRKBGtxSMdOwqayszAa4ACQ+DT0Cwl6kMEZlIxS/WpJ8eJKKEpkimC1CDtke/rY6lL6Pc0umdzPHJyA9465LqABcGH6D8Uzy1EkgIEwZMipS4Tkre42n0JwL3tp6SNC4lMhUtXlvO/Xgb3Xb1Op5sVXQRkMFkHAJmywmHu9V7Wy9Te4N27/+m7Xv/f/sqvvfec2oU/9eaXU6HxzL2rxY+LyAuzLFuFUpDMIFMGtgpXHji8dHXO9qbjDz36f7/7La/6wN/8rT940m+cWhBKcfn+y1VVllc5FZ6vmVdmM5rZPhCAifhmEzyjK0ATywKVsh4GC1B7P5W2CT7qpBGA4GCtg9EaCNNsgSclKoaIBc/4FSEImDwUYgnMkAJRbOxrDsi0Ql500O/1sNwtkLMgZyDPdNS3UwZ5YVDkBfLMoNvrQnPyQEopEhNDswIrJNr2DINP5kVMZUa2ZwpEyUQPYaKgvZ3VN2tbTlgs5hrLg4CKfL5pCZKRwHp7WTKgGYAlEhSGILXFaidHZgy0yeB9gJwdYORdBDVmuAD4EId3kZxfoRjEZrWu6xfC2Y9edeCiU19+7MF2iLWN82RBr1nuF/SymvCcXqa6TAGsNZgzgA18XaGTGyjKu5u2vK7Tzd41HI7vB3DbuXfJ7nLv3Q8FpZ9XaFrNGVC5BvICVgATAHh/pLu21F8Zb5pw0g8AfKQFoW+RsM5eZtn/oCnyK5iZIjWZoVTSgqNoqhblYVJNa7IAMihqx0x+NrHkEcCTwCVoConSLCIwSiH64BDEu9gQSSTi2LOJGQaLhxGBIYIyCtqoyELTGkVmoDlK2xRZhk6eoyhyZJlGr9NDv1Og3++iyDSMNlBaQxGBGVDaIDcRLBUkOb9O4UUBO+wjZg3pZt1eZcbGYZbhFhWyz5fKp3omEcjv/F1jh9E8z6xSxJxm3SyIEYHSAC4TUGiG0RkIBmIBVzuc2BxHqUDWUdaHp75QksgSACDGHHVcvZWt+8y1Ry75zB0P3yftJ6aNXbMgosuW1ldfC60PaZ2DdQbWGYRUvKIUAR7IDCPLi1U22ZXF5vjqc4HQz7ztVXvhy1f19hx4BZlsb1AaQamJK7Nmhs4VXF1BRK8Ue/bctJf123/hLbfc+b/91h+ebEHoSR5XHLzyYOnKt7PRL1fG7GsW1sYFNaoGpDmYpB7AzfonaRcfOMrEpP5NM1MjFJvpQgziSDmOap0erqwAseDmuBKlOhUBigjG6Ag0pNHVjF4nx1K3h36/H8tpnRzdIke3KJDlBoXJUeRZZLk1YJastZvXQ4woQR1X8aTLlhzAJcTyIZo6W6OwwDvqwhes1kAT2VMA55qdmhdCnfw8NCXARgx2XoOPmOZ0+WYBSdJjjFIQT7AuYMUo6P170j1P4MSoxMjXUMRgNghCCC7+jZqyI5HqcFHcVA+Hb9XOHAfwaPupaWNhFvS9rzuYGbwqkHl6rjSrrAAbA1IaLkRmp9GxNB+sBQfBeDjuOOvWfuZNLzM//p4/tjuO+f2vyfrd/Lmms/aObr9/KTGBjYYq8sn6lBkDEkHwjFBZCGGv7hRXFZm5BEALQk/muOrw1R3r6ufC0Bu1MUebRayxY1CkEJIYJzjt6YUgkvhcSVcuBGCS/hAQKLK3fCoNhZCUuL2HkijOKcGCxKGbGRgDGGhkipHnOfr9LlZXl7G6soK1bhereYYskQOUUhEEmWIPh+KePYpFyySbidkZEFLzhijZaTcImtBSqei905TOpiZ6U9AINAWeiVPrzNzOHFlk9p+S3FRJUv9n8YBtk1HGbKTJMtNzCkNIJiZ5c+W8VDojmXWobXYBM75FIlDeQ0NBmwyyZwVOHPzjpyHDcZyRIgWSqA6BRL33wcWSrMn2S2FfG7z78LVHLjlzx8P3td5DbcyDxVtft7LeMa8rljpvAXCwU3SgdQYoA1EKRCFqI4YoVVWOR6hrh3IwknJcVta6hVYiRuFYr9/9S7roPT3X0RqGjQG0BlhBEScZrQrWl4A4uMplvqr35EYfAfCpFoSexFHX1bGa3Nu1yS4DkZ6W4aI5HVI5KdpFNyy1OGcSyQQK1BjeOYA4Ga4lAwJBlK9RwUVH0NpCcUDX5Mi6OXqmg/XVZVx67Cg6mcFSr4uiyGFUU4IiZMQoOJqzccqoGvbbVDonle+8AKzAisCKJky4IFGxOmYPSGrTSbTUpwV+RsSUELOMiWU37cxkKCHZfItsOi81sbKgbcgEmTlWmAOiyfAvI5U5tz8nTwgIc1nZXJ+JmrnT+DpdfF8UEyQEwJboacLBtSXUwcFLgNsaoQwWQPQeAhQC3ETVm5iIjDnqxb7JO/8FAPe3y24bTfzkm15NSx19ea+fv8H0e9eSOBRZFs0VualGKIi1sOUYoa5RjkfYGNVwVT0Yl/WJv/d7H9xBInj3225Z6hr6LtLqmZmijmGCyXOwNnBBoFTsHddlCSc1BqMB7LjG1sYA7DwF5570HllPaRC68uCVe8Z29HoYfm4QWSJM7RlU2gmHVK6aNNnTUhjngrZVniSWukR8aqMnzTTxYGuRZwpaASv9Do4cPIT966tY7y9hZamDXqbBJNCKoNLiyUwgzeCoj5Pgr1n8I5hwUvAmtS3DoOgjJD6AOZbdFCfYkKk7aRPMBGKdymcRVhmxtxUmPj/zRTWeq7rNeiNN7bojb3zyLNN+2pz3Q1hcxiMCBdoBQrFPNA9esrASGEkhpBgSfCx5siBYCwXGcsfgwOoSqqpGWdXwZaKMKwUfCAjzfShitSo6fKer3LOuOXTxiTsfvX/cLr9tAECmaKWX85s94XojvpMXedwwkQLrHMHHmbzgPcRbjMdD1HWN4WhoRxtbxwej+qFFxy00buz2Om/P8/zSItdgpaJ0WFaAKR5fQoAXh7ouYW2F4XCE8WhsVW1PV1ujJ73s1FMWhK4+eg3VVXmNaHqLMuZoo37Q9IFAlHo6zdIXhyQFASFhQki2bSE1sTkIGB4kHhIcWAI0Rcpwv2DsXeljqd/FSq+LQ3vXsb6yjG6WoZMZcPCg5K+jktcPhCDOx50U6bhi89TaYCrAKZOlHxPpGwaxillDcCkjUVMUoflsRtIMkSRBUo+QZnxkYqJ0IWKpsyrdOzInmpxlBDqRif9SY7knErYZ9PFOkJo8bqr4gKZ/k45DIHCIZdCGKOJDNLiLfTEHDYXlTGNPv4utUYlxOYZA4BRFBl3T76OZ16PUkSqUryPLt6IVOG2jWUjJX2FD/Wyj80MCB533AcVgbaCUhncB4izIWTjvUVYVKudQ1uWp4WD4URvUA9uP+Ytvu2V/v5u9hvPiJsUCpZqPcIBCvN6D9/DewTmHwWgLtS1R2Rre1mdlVH5lOBo90ILQkzScswdEyZvAdBkAmlg1KAaYIn26YcAlwzVBmg8CkiVALGm5EE3ZNAQG0bqAnYVhwkq3i+V+B4fX+7j48D4c2LcfhYo7dMMKmgEFm7KKAJKYtUwWP6JU2AOIUymu6c0QAyqZ1s1aPaQLVFJOExk00b10to/SQAYrHQEXlHx/KJXgplnNIsVvSc9HC0Cp8VgSCRNF7glEpeNOH8loUjTBvKZe7P80g8FTijwRTwCrISg0PbqYJEUfJaao8yfEgCY4HxCIQIrAEpCRYM9SH14UBqPjqIYOpDxYKQTi1OydOrEGyIoofq4Eee7VBy8+8aXj94/aJfipHT/9va9e3bPWfTNydYXOdKYyHRlwRseNqos6iyEIgvMYbG6htg5ntrZCORx90Tl88Gf+8KOntx+3k5ur9+zd/+KRhD25UWCjoE0OY7JoqeLjZ8Y5h6qqYK3FcDTCuLSh3Nq6n8b+oy6EB1sQelJmQVerqhpdZ1V4KSmzJ9b8OdKvsXO331CrU0cCLkTnTx8EwgBJgBIBgoUEB42ApY7BnpUlHN57APvX+rho/wp6hYbWAAUHxQRNEmeGJNKl0cyocFKoJkRWHRpSQZhkLhGEplkMEnA1THFqvOwCQcBplokm5bYJtbmBAyY0pOTkeddwLtLVvjga5YVFHkmTAhrzpJRH1JT1ElFD5gFs1pm2mROaOtbOlvFoQgGfABFhjmI9gdoEyEEA4fhv8VHdIWNCL9PYs6xxZJ/DOJzBmdpBKQazigAUtr1iow/a2r+Cvf842t5QW4pTuBwKN1JmDud5Dp1rkNYQ4rhGiId4D6krjEcDWOewOSixuTk4Nd7Y+rAL2Ze2H/Pn33rLwW5mXlV6XF50cmgTiVKsVRwaR6yTO+9grUVV13C1g609RsPh46GqP1yW9gM/+YFP+Sf7+/eUBCHn7EEP/1bS+uLpQsbJ/jlZPidZnskCmSjEgghALviJ8nJ0Bg2Ar5ERsH9lCRcf2Idjhw5g7/Iq+rlCpj0UB8BVcXFXKipR62gzLZQGXongOe7UQSoqXifMYGoW5lgmbCR7GuBpFmeeDFxOM6RGBSBmSmoi3Nmw6oQWQQsADjv6MgsLcGkuZztTjpqsanu5bsZnaQ74ZQJrE6CaB6FZejmlkuiMHcZs6TBRu2mSxSQJIGE0eSIBMCLoacaBPWs4U9UYnxqgRLQFF6aktj2VHFI6XxFfPSs4f901hy45fuejrZzPUzX+wZtftbS+0nuV6hTXdrvdPO/kUJlGlhXQOppeBuvg6wp2XGE8GmM8LrE5HIXNs1v31cPqg7/8sdsenz3mz731Flrq5s/ur+/5blFqr1EGWZaBEtWb0m7LBw9X17BlibIsMR6V2NoaOrLu9vGo/q1/8IFbH/xWeA+fciB09dGrdW3Lq8Xw80FqNdoyLPD1mWRAIYlNhyQbIwjeR6kcilkNU4AOHr1c48DqEi4+sB8XH9qPfctLyJkBcVDJu4e4KR8lnx8QWBkE4bS7j+VAIY55ycxAJmha/pIZETieLMDT3kpDoIu21yqtzc0CHe/XLNhC0z7NHA7N/2MbsOz4YaSfLijNYVpBhEyelmYyrlngmrXwns1ypnQIER8hqiFRTPWN5lUZSCazQs3fMz5eIsGBAnwIEzBa6his9zvYGIxANqAMMcsMidIuYeY8tTrsQ7jFeX87gEfa5fipGZr8ZTpXzxNSB+Ncn4HSsWSmlInbLfGo6wp1PUJtLTaHI1S13TCsvxA03b+zuuAvFYSXV+BrO1pDZxlMVgCKIaQgAjjxsNbC2hq2quGqCt4F+LI6IVvlx12Qz3+rvIf8VLtoQnB7AoXXkNKH46LFkRlG21Wxk2CBxEXSC2AFSadMYAjQwYNtjczWWC8Mju1dxdVHD+GyQ/uwp1cgEwsVKmhqWHJRZDTK4GgIGF4IPs2zCKloPU3ReE3Q1NQ4ZQKcsg4GSWLNEaNR++bEHOMmk0kVLybMgOzUQ4co3ZIOHU3mcDD99xwQzMv3zA2NJlCY7U2d26wv9XV2ZGEXEoSdtIfZ8uLM62VJYIRE/KBIc8d0pog4yiBp9lguDFazDIU4KIrSP2heF830w4jXguLnO+8vu+rQxapdjp968fff+PLl5a5+tRO5OstNoZWG1hm0yqCSOoL4OJgu4uCCw7AaYWQtqtH4ITd2fwLw3AbmZ97y8rzXy16me70XQqvVvNOBzgowKSjSsWoiAhs8nKthbQ1na4TaohyOnBrXXxgPxv/lZ//0098y8lJPuUxIgj/mKTyfSK9xYsBR00CR6SI2GYuhCEYhLZqRmSUg7yG2RgbBWqfANRdfhP2rKziw2sdy1yCjOJSqiKBIxWwEDAlxh66iKBsg0VwtMQ7if9L0gThCCk0bPcQ8XWSbXgvxREt7ttfTrP+KuJnGmfxsjqnGlNozTUYYUoYSZYWCYGE2NDvbM/k38ITM+mYMJnYp9U11whdlWE3PKW0x4H2yjUjeR4HDTH8oyiuRpAHeNMxrvUukDcZKt8B6v8BgOMI4EJxiMMeBXhemc19ExMJ82MO9KPhwJ57kU+ltfP1DSX1Fp7/0IjbZoU6eQSuFXGdQKoNiFecLxSMEhzi2HuAhkOBOudHoIyHgY7/4kU/NlXK1kks6ney79erKFUXRgcmK5MOlQYrg4OG9h/MWpatQ1xVsVaIuS1BVnSygvrIJuudbKpt8Kl00Vx2+cql2o++A4WNERMwM6yxIR5Zao0w9K9ApIbHigIlUDwUPCg5aAvb0u7jq2CFcefQIlosMnYyQsQcHB8Upd/FIOxkD0pyGXxFXQmIo1pE2kDIcoma3HhdNaVhwIEiz4ApFYOFklSDbMxOa7P7BnKjjEQBjKUpmvk/ASJSGVuP6zGmYVRaM8SyyKA8i22wm5utwAixQTEhZqMwCqMxgEs2VBJu+3IRXxyppyUXiBROnjQXQ9I+IJMkRzVPEo3J3HCJWzPASUGQaq70co+UeqkGNWgCtGAiMoAg+8ET2yAvWIf75maffaUHoqRU/9eZX7Otl/rWe+WlFpjuKgCzLwKzAaKoScVTDuRpVVaKsS1S29uXW8C5v5XeJ9Zwq+y99/6tWlnv8es6yZxute9poKKOhk+YjEDlLCBbeWdS2QlWXsFWFuqxrPy7vGpwdfvCnPnz76RaEnqThnNtjg3uJNv09RDxdjiZD/QKGNEppsQQj014DiYCDg3YWOXv0coXLDq7jiosOYq3QyJSHktgbaXo7SM8TEiNMJc/skJhujb1Bw+4iYNL/oMRcbr7KBGyms0LzpbEZGRueyR4QtesUKQh5UFAIFCJnjgKUKAh7iKiofyfxfiIJ8Eh2FMO2K2JvB51mdqexbQA1KgbSTARN6O9IlhiYlATDNA9K4NFoY1PqgzU9ofkyIyJIhwAwx9Kn+DhvNTlfiXNePh4zUtI1lBA0BCQeyzkjrHax5TyGYwtiFf2QlJp4GMXn5QLMVwBy09UHjt3/pcceGLbL81MjeoV6+ur60kuh9MFca+QmB1MGojjwLT4gwMMFh7IuMayGKKsKtqwf59p/VMCfe/eH/nzug7W83H3B2p7+91TgyzqKkKkArQikFTxxmnNjKCbAxjGQUFco6xKj8ehxqfzHx04+tOh8/9EPvCHvdrID/U62P8/0Moegy6ra2hqWj4wq/8D/8h/+i7Qg9E0IIjkKpa4g4gwUBxKZFRRopieCCfDIpPdAaYhUoCkgUwF9Tbho7yquPHYAe/sFDMW+AqUFL5Ca9HUmMzMk8DQzjElNnypEtlyz4KcFO/rxTEGJEVKJDkkxIKk9J7JDI8ND20AjJE+jkJhqgak5GkBq+vNkQTH5fsc8zyQN2uX9nYKOJAbPFIAbWAkpC5uz+Jv815AIZoqKKRdiTG0aUglSQqLOT5E6+gElBQVSUJKaw+QBjucSQojvQWgEXQEJUbwVEtBRgMsZ/UKhqCwqBIgiaDBq+LRNSbNjpNaDc89x4t8PoAWhp0Iv6C2v2FcUuMWTXNHRSmVaIzMFWBmw0pF05AHnPWpXY1yNMCpHKMfOb548+SU7qN/78x/6zJwI7i9+/6v3LS113z62uKZXZNw1BpmKElVQBEexIiLBI1gHVBVQl7DjEcrReFiNRreNB9Vv/sxHP/vY9vP9x+98096D+9fftrzSeWVemIOGuCveM/kwOnXm7MOPP37m1/7RO17/wf/l37/3ZAtC38C44tDl/SD2BpDaNztfAjSzI8lVEwKFEA1rGv5yAOAiJVuRRyfTWOlkOHbkAPaurkJRUjsgmaEK80wpiSZ9psl6LNPMhbYt5M2uHgtUpZEsF2b7MZj14qHFbDYCpyyKJ5oCYJordIFpR5msoYjv3pPBjrKczCg4zGc2DSJJwprpQJLIlGwQnWppSloIiFYLk6UfUeg0RLXwhjwSZsBMmhmkyazRjJRQIyuEOIclLLGBnACOmZAZjaVeD/nYw9cOngieAMUM56dUdM9YdsDTtQ970aprPyUi03S1LrJnAbRXJZUVH4DcmLg5TNetDwG2qmFrC1tZ2KraRF1/xku4a/sx84yvVUZf4knvMZmJ0mHaTNRbmvXJ1RZ1OQZB4HxA7ZyHhPvFhvcHVndsP+4vfN/r1tZXe+/Iuvk7qiy/QSkumoF2YYJZ33P1itL7i2F98B+/8y2//tf/3W+dbUHoGxTeu34gf5Mypi8zPR/iNG1PzQY8Tein72PPJElmOIciJ+xbW8bBlT72rK9Ba4ZYC9Kz2mmLiM07lu7JYCYatYbZ+RpEdYQISLRjGHTnLA52ldeZZBMLgGpHOW32UU8gQV+kjt0Ek8wlT/N3oxlImCoohLmsCkkqKZEKkqq5NJJ6DZURM7ekWj5b3mz6Q5NxonRe0njrhbQpUNGdttvVyM0I49JOthNKMZy46ZSRwDimIzrghsv3XnTX3ScfbPXkvo3jx9/w8rXM4LurQFcsdzuZMiYa1imNEHycfxNCCBQp1GUNV1r42sGV45PwuI2UmpsL+qXvu2X/6nLnnWNrryh6OdjEYVdiNVXqD5Hg4G0NCR7WW4ytR+3cCTcqP1R5+f2f/dCn59Q73v2213RWl7tvyIv87arTeXamGJlWUCrSvENgKBV6elXdTNmYu1W4B8Dvf7Pf06cMRTsEv+4QribF3dlyGE0mNSM1WojghRAkZUshZh+GAjI4rPW7OHpwL44d2Y9ekUWFBMVgwsQEbU7iZhu7aztwzMreTDOhGWmdbcDSyAvNLuLnB4j5cyLZCTALQW2X759wGVQa1t/CqaOZ0mdz43Sb+ZnMvI9zYI1JsY7ToC6TQFE0AqfJsCnN9M1k2v+T6EjLSRKpsQ5nBjpGo5dpaAJUU65V01kr4ZgdCdGKR7gqBN9pl+lv7+gYXGfy7IXKFAczk0NnOZTOoU3qGyLAOYvK1ijLMcrhCNWwQjUYbdYbg8/Xzn/qZz9425xnUGboad1+9yZSan+mzSQDIqWgVCq/BwdfjRFsCWtLDEYjVFU5QG1vqy3eE1h/ZfaYP/n6l6tuYV7ZX+79CHeLZ3Y1o5dFfzKdGeg8A2cGxhgUJjfdpeVL9u1bf9M/f9fbDrQg9A2Iqy66ipXii8F0kJl4Zos+Yx8gSaMs7cwbejFRtLy2JbpacGBtGXvXlrC61IEiDwQXyz0iO2wHzgVCO+4nO20SaJt9woWAwRMBDFqQOdG2OZ+vFoh2vJ5tzLnJvI1MgSjIdjCaLWgmu3OZ6Gin/zgN68YPqwJjwk9qNOVo0W2qpkCYH4qNJb6ATDNWul0UhqGbjEoSfZ0iwEExAlPPBnd58C0IfTvH333Di9eXe+ZNed69ppsXxrsAxTETcomGHXyAdRZVOUJZjlCOSlTjsR1vDO6vh9X7AniuFPcLb7vlSL/X/d5RVV/d6+TQWWTEKa2hlE6M2YDgLLyt4WyF0WiEra1RKMfjB8pB9Qe1D5/8mT/+xByHNdf09H6v82Oi1bP6hVGZBnKjYdIxQSqqgTAhY4ZmXis62RW93FzSluO+IaW40CVFVxKbFSGFRiFOI0m/pN6BzKklTPfojABNAftXl3Bk/xpWuwUyTiZpHKIlNfNUImdCEabdMw3BgmFOSj0Y2jXB2a7Ptv0YOwzmdgGIyPZL39PuQPO1gs+sp9CsCd7s/WTyfs8SEuJXTgy6hoAQUnmCU6YazQV9NL6TyKaLLaeoAB7Ep79LQ7KYZoLRmyikyt1ERS8qogPQBKz2Ojhd5CjtEMoJSEKkxUvDbmQIS+4kXKTFrQJ4uF2uv/3ib7/2u3VHh2drlmcx08FunkMEyIsutDEIwUY5L+dQ1SWqskRVDjEuxyhHw9N2WP6xDfwHP/+R2+fmgjqFvrm/snKzFdvXTFAm2jWAdVSx9wHOOthyDFuOUY5HGI5KVHW16Qfj28aVff9P/tGfb8we8+ff+uqre4X+H73Rz+l0TF5kKjqvNisf6SSKHBW4UVs453QoyzzXarnNhL4hIOQLL3IFKdVtSjM8ufGcF440hmgiUJRKNRBkDOxZ7mKlk6GjCOSiVUMzvBop3dPsZ/t8y4VnLxf+uG2VqW9YnAuIdvvdFGgiyIcEJLIIoGYoBw2RIerxSZQ7CgLVqD8I5vKjSGpQUfYIGoGmN4FO2vfNVzURPm2IF5yo9yRhxuKIoInA4tHJVMqEJInAejBHEA+QyNIj6EDYLxKOXbnvsG6X7G+/UCRr/UK9rtPvX9UtjDHGoN9fArOOPpLMcN7COwdX2STTM8aoHIatwfCE9/g4WM9puf3S999yhUJ45aiurjW5AWdNKS5LYwHRhNG7mAHZukJVlajqGtWofKwc1R/wwnfPHvNnvvc1Rb9XvK6ztvbKbq+72imKWFHQKasiA4KGeMB7j+BqhFBFmwlf23o8qttM6BsQzrmOh70oL/J8MqxI2+yh0y5bJDKgFEWhUhUcFDyWOwZ7V5fRyzQoWDAFMAI4sWBINZpkM+6emFeZjpP9DBFKCtjTctTitZwmLD2ieQWC5ng0T13b5jCKGadR2bXUdj6gOZfywez5zN5v4pCKlCWGMPEsYsLE3oEp2mMAkSQiQRCCQ9NhkzBjfkcUyQOgRPUGvDQ2FbNWG5zYcZKAx8EHn4Z0dRxADn46u5TYhSo9HyXHWu0FGQIKRVAUYBRBBRWHVYOASM3S0ldJ87Ui8mEAg3bZ/jbKgl73YtYor2fTv0Hn2YFOlqOT5TBFF8QKSkfXY+csrPUYj2s4X2FYDmDr8SZ5d6sn3PYPP/SZiaL1z33vy/ctd/Mf4My8SiBLJu+ATR4VsmecgqNXUA1blRiPR6hqi/Go3JLafa6s/Sd/6k9uncus8oyv7Hbzl+pOfrRTZGCtoIocgRQ0GzA0rA2QIIkM61FXY/jaDeuzZx8ZDgaPtSD0DQjxvhu07IPibJo9UPTkmChL0wwdOUwYVIriRM36yjLWl3rIOFkxJCfT2ZKWTLoXzfx+44S6HVgwN0x6njxkrkS1qNx1PgChRvngHAy7WfA4X4ntiWRpIUzfl9BkG83xggCKk71DmitKgrHUDLUywyc6d0gSRUEA19hrKIL3AusdaicT4CPipFbhk+RJMswLDuAw8W+S4CIAJYAMxLEnFAQsAUoIy90CuWZsDS3ERzo3kZ6nySvV8yFc6X0oWhD62uNf/vffrxQTfuRf/MZfuBWBVnRwdan/xt7yypWZUmSMgdFZuq4iCCENkvo6IDiH0WiMsqp9WY7uEx8+DmXmMpa15d7LOr38JWyyS1WmQVkGlUc31mYzF5yDtRWqqkJZjlHZGlujsXXWPSxW/lyg75vvL71mfSmjV3CmbywyA9PJAK1AJkMICi4wjIpaDuJq2FDDVTW8r0HeHq/H5afLunqoBaFvTHSVUr0gyeJ6onGGGRtpTJrb4qM+U0YCwwE6BOxdXcZytwCHANUMWwYHKD2jXZYWW5qtczZwpL6G6qdsmwuaz1CmSj6UyoPbAScVCRdQvRt8a9xHLxRwzne/aWaEKRynQVGZyPTEgeEQ/JSuDgK0SWXUAGgdzcCSzXgAobIOg3GNcVlhOBqhth51XaOqXaTJioChYRjo5Rr9Ike3U0ArFTNgNhEcg6QBwMZDSaLdRogFQZ2ytOVeB/0ix+lhCSWR/ACS5CuVyOWsC+uqSxh+Da2EzxOOn3/H9+lMyVphcGhtqXNpJ1P7NTP+69/+y2MBb9YuPD4Y1w9XTk7/d//i33zTQP5/f91Ls44JzyqW+s8X1ocykyMzGZSJUjqkkiJ+QMpcPMrKoqodxoPxyVBWH6gcve/dH/7M5APz7u971UVL3e7bRYUbMgZUbsDaIAQGm5hVBS9w1qEqS5Tj2FsaVhUGW8MzUtoPD0f17//U+z+1Ncms3vJKXunnb1pe7b9LdfuH8kJD6QyiFIQ1oDR85RGcg0hyY60rlFWF4XAkNNi6azgqP/o3/vP7By0IfQOCmbqBVRFXv0gg4DRcKjNU6Eb/jCmxucRDg7DUybDU70ApArydettMFA9SSYcxAaALIQgsXry/GoDCxGMEi+R0tmVCi7IemXosPGHg2V6KmwcgmZm/at7qWC4LEhlmwmrSM/LeJzfWgLKyODs8jXFVYTSuMBiPMC5rDMsSw0GJcVXCZDm8D3DOR0Cb6UVpCHrGYLnbwfr6CtaWeugVOTqZBitMM7PEHZcgM6SU2BOkEJArjaVOjqUiRzW28MwY1tHsjhr9BOZMiI56549cvu/w3Xc//khooeXC4ufe/rb9q/38O4uCXtvpd67vd/K9mdEdxZq8d5aJyp5goxgMH6pH9e3/4a/+6Ec3RtXnfuz/9+8e/0afW85ybKnfeTvp7OpOXqDICqg8hzIGrFI5P8Tsp7YW1tWo6wpVXZd+XN3pav7P7/7wFyYacT/5xperlZWlN3iSq7tZvppnDF0UUFkPPsQB6yCC4C1sHYkIg9EQw/EYm8NxVZXl3W5Qv9cLzw2m9nr5Tf2V7g/obu/pRWEiYSLPEbQCkYbzHloxvLUIEhAkwHuHqqoxGm4dt6fOfGo0Dl/8C8k0v90v8EsPXMre2yUQZfMDkVO1bE61NxcklmGYoQNBiSBThP3ra+jnGcS62MiegAwDrBC8T7OOUYB0orbQ7O0F5+caSCrczfjmTNx2ZKfF9hQUaNovOk8mtL0HtAOMgkwyot2AR2Qqq7NbP2iO+RbrcXGENIQJ0NkQUDsH6z1q61DWFsNxNPyqrUNV1hiVY2yVFaq6wriqUNUONgh8CMlTJcAN6hn176l6RMxUBcNxjTODEU4PhljuFVjt97B/zwrWljrQSkPg0LASo74cJ928pmcVLdc7nQxL/QKnxhWUcNQHDDTh3AUBAmHdS3iGiNwKYKuFl/PH33/zG/eu9rN37D28/k5ofZkmWYnZRez7BUhcnJUCL/VvzHvynVltX+1d+Uf/6kff8Sdj6z/zV//tf/yG2Bb8+Gtforvsnt/pdZ+pjennJofKCmidTRxOQwgxa3EOtqxQ1WO44DEajk4HKx93QX1h7nOncNHK6vJrA9yxrGOQdwqYTh8BGkWh4aoysuysRVmWKMcjlOMhBuMhhsPxWZT1x2ofPvfzH5w6pv7sW16x2uua7+csv0Zrji6seQalDTRrQADvPDwCPAV4ZzEeD7G1NcJwVI3c1ugT1uK//R9/8PEzLQh9YzpCioj6AtHzQ6Qy40ojSf0W0YCOEjMueLAA/U6BzJi5xVvETyaPo84aT7s3CQAYmFgkPPGciC4gG1mg6bYgE5oFsJ2/2wlMcs7n3Umv3i0rkjDjWySNZXm0PB6Ox9jcGuHUxia2RmOMK4vhuMSorFE7hyCCylrU1kYjwQB4EYRA8CD41DtinSeNOkm9PJ70nYQA0YQqOPhRhWFZYmMwQO0tiPdiuVtAE4OUjjjkUnltUqYMkQkXPLpGI89ykPcIAVASouCrzHguKV4mHW4MIfRbELqAUtdrX607Ob+4t6f/Lkt4Rp8EmgR5ksJRSqEAooOo8/ASCq/o8IhxaPnooUtx8vR30ebw//lnP/R97/+f/9//+HWXTDIcDhc5v4SBA0udDrIsLuyidNKHjPNkEhy8jTbbSdm6dmV9dzX27/2FD392kq39X298Wb7UzV5U+/rSrNC5LnKovAOQRjR6YTAxnK/hXQ1vK9S2xLgaYzweu7oc3Y8q/PHPf/CzD8yeZ5Gr55Gi52XdzoFutwPd6QKsEQJBI/a1wYyyHkNEULoSW6MhxnUNVKMvhEr+07jyn/kL67l920NQHCTpCkT7hmzQLJYz/jogxH5Rsn5uFmUCYLSC0VOL59lF3Yck8Dmx075gYvY5S3K0IH3aTa5narS2OBPitCgHWpwB7QCk7d/SPODQ9mxn2/zPpLEKH+0gJiDBqcxW4eSZs3jksRN46JET2ByWKL3ACUUSQgKGqFbCsXwQZgCC4i4UiiJRQJLWHLix/Yv1eSHUEsCsY4kDDlLXOHV2A53cgElQGIOMJVH1o7utcNQLJAbIeihiGGPQyTJ0iy7GwzINzs7IHYkAxF3S+vIQwhpaHbnzL/IK+/rL2fdkneKqQhE6KqDICwTOUAsQKEDHQcro5+RqeBFIpqiWcKCzd3VJ97K13tAe/uUfeNOv/LVff8/XTUD2b3/Py6mbyzOXVrvXK+YlTQStDEgZkDYgxXEGLcQ+ZG1rlGWJ2o4xGm6cocp/2gfcN1fay+iqpbX+O72Sy1kJTJGDshwMjY4pYJ2DIob4EDOrZFpXVxWq0ehsGJWf9D778lwv7a23XLW83PtLptt9hkiARWwnKM3QUNCIsmIQC2ZBZSvUrkRAALv6/npj9L6tUf3Bv/tHfzZoQegbh0IMkpxJsUpzJoTpwiiSVpsQICE2nQkExQG5BroFo5cbGGJQiLtyZoLiaEbnnIfW2URpusGO7RQE2mVhb8QOm/49T1AgLPzzbBcK5SRmuuOJmqlMiXYNkyOLn5uLauyuF0eYlAqnJbrFmdCOAVQkVQPvkytgQCAFJ4JhWeHk6bO476FHcWZriMoJrCiQNgggeE8Q72babpEOzdxQoj18EIgPUEmqRxMj1xzp9ekE6uBRNjTx4EEIqL3FybMVgq8B8TiwZw3QjIwbEw+avC/UvFYJ0EQojMb6yhK2yhrjuk7SQmoy/0RQrBSti7f7rtx/WH3lxCO+hZrdo5uZff1+75K6qrrrqz0oiQu6U4A2OVgRKGUaEA/FORgeAdGry5W2q3u9603h33XA2fEvv+11v/bXfvP3vi6lOcXYm2XyndDZxUu9DrTWyIyBMhqkdJwUCIh2DdbCVakXNBptcu1uq0r3eyAzyYJ+5q2vvLjI5I2BcFNHMXd7SwhkAEQjPBZBroFx5aIHkbWwdY26digrP5LK3eqdeo8oNQG2n3rjS/euLvV+wBTd7+gWnc5Sdwm6k4O0mTJwJcD7GooEcDaW9yJzrxqcOH7r1unh7/zE+z7xF7phegpkQiAQshACc5pNIVIQ0nBhqn6tCNDEkWRAQCCBh0c3K1AQQQU70SWbZBABcXdEHPsDSfYlzgCFSXbCiRSAEH8nmhGEUmYSNdKYZWLmpiieY6PaE9lXs+U0BlG0fvDep3JiUkCYIQREgItaeJQsK0ABmqIvTrSK0BGIGl4DJ+wSD0aIHzaR3YxPE+415gaRBg2Jg6YiIdqa+xAf7j28AOO6xpnBECPrUQVCKZGNRn6qdM2ILrIKSbA0OITG5gJxRkslGZ2O0ejmBof370O/00Uvz2OZTRMCC8blGIPhEGfOnMHW1ia2trawNRjgoeOA9w771tex1Cni8DLr5ERbQ5zAaAXvAliApa7BisshxysoDdQ+QEjFzM0DcB7B+eWc1TUScCtaqva5awFBjFQOvV4P3jkQWagsg9IEVpxYpyr6WoUAgQcFgYGFdQ7LHYPKejOq7VWmo95RKH/PL7z+5X/4v733fV8z+Hcyfnp3pfc8zvReUgyVR7ozJ1o2EUBK4EqP8XiAcTnA1nATg8HgwdOPnfnXwsXHfukjt3kA+PtvfEVvqdBvKPr527pGry8VBTKdw2TdmFVBAFTwrkawJcTVCN7DO2BraF05rD9fjfHPAmcf/Ucfui0AwE+8+oW9boY35R3zZp11Lu4Uy8izLgwrCBk4AjyFuAE1hLIuEWwFPxyChVGePP0Vdni/F/ncX/R18FToCREEKg6iBMSRxKnRQHQ0jT2eZrGPgpsMrTQ6xiBP3PqpO2gSbU5WBzgPsUwoWmw3IDJp0KcHBXhQSKIaHOeXpioMO4dKeXbGiKaMv6gKHSaK1NTYH3C0bwjBA8FDVIDmpJPnLYQUwGpGvGBK7GIBwi7Z2LR3IruW5HzkQidfoZhlGGXQLbpYWlqGpxFQ1qj8dL4HImkgNNoYMytopcAMGKWRFxq9boFOJ8dKr4NenmG510U3N8gEUEpF0VHFsLAoa4WwvoTq0F5YF3Dy9GmcePxxDLYGOHXmLLRS0JrRMwagWAoR70ESbb3JOyA4sBAKHTPjzdEARBlEhTl9QNFm2Vv7jBDCe1sQOneMh6PNrTN8ukZwaq2rO12FuiqhkcHDAjCxNEoc58lC9MzSJm7iSABwgNc681l+TabwTg13P4AvfC3n9Xde//J9mt3LoLMr89wg72ToFAVUlkfySgiRxGQt6qqK4wHlGHU5OuvH9sPE2Z//4kdun6ip9/u961bWOm+sQ31Zr8iR5zm0zqFUnnq4Dk4sgq8RfA1rK9TjMYbjEsH6E35kf8uR/tgvf/i2iZpBv6dftrzS/+G8U1y3uryEbqcXCROsIERQ4mFDZJp6W8GWJWBrQAiDM5tb1cbZ20aD6n1//4/nh11bEPqGYNAEOqYlqW0lpTQkkno7UyuGzBgUeQalef6A5yQaNEs2z3xPqT8SjeRYGJSkXxQBJAytVGpyTjhBIOYo5y4hycQnX5GJ3A0mXjqNbJCg8TJqtNYESlHUo0IASVR4AClQCFNWXSp5ScC0rwKZa18tYsPRwr5Q8vgRSQSC9B6IQIRRKI09/SUEF2CE0GGNyjrUIcAFh7quIVqjMBly04NJAMRM6OYF1lf72LO6gn6vQMfEeaBunkWgQICCwDsLIIC9wOQ5QEDtM1gv0MzoFjlOnjyJ4eYWRsMhBpqhl3vIlAIxQ+sc7D2qcQn4gEJnsFVAVxkcO3gYo/GD2CwDXLpmHANeMQJkWRhXay9rAI63ULN7lNadLkt7l9vaerzT4UNsskizpxqaCIp4TlaLkveTIoqkIB8ik5UAp81qd++eG4nPvOiX3vjye//G77xv9NWc0//+mpdRRuG6vNv9TmOK/YU2UKzjoLQXKJMqGyGgrMaoawtbewzGY9Tj+vjg7PB3f+Ejd0xKZv/gza/qLS11Xs4mu6hHqsi1gtEGSilw2jwGUoBXqJ1gMK5RlhWqSEZAqKu7faCP/fJHbptYdv/kG1582ep6/12617u20+2h6PZgJcS1REWgDiFKXomPpAlfewy3hhiWlfPj4ReWOv1bqzLc/WS4Dp4Kc0IiMhF/mempzO/sgwiYm9Z2XEyV0jB5BiKBExdLcdvJAhfIfIuUXwYrTGwNONmOkgisdVCaoZSJLqvM8AR4ifRvrXQU5+SYpQkSpRicBiYJTiRqTUlIro4uNTuBPNPo5BrdLI8Xpo+lDaViT4NCcj1lmoCPJO0HWdAHmgWkpj8VQlNOw+T7xoJBGq01H5AzYW2pCwVAe49NrTCqHUpvUTlGZRjaGHS7XTAYhhWMJuTaYKXfw561VSx3C2QqKpwTBFSPoTiVA7lRyCYUOoPzAd4JTLJTp04XmhRQC9gJnK0xriyWAkBaISCgqutIu1cGEhhEGoo9uPbIRcDOQ0FSlqchTGnnCXLEh3LgyOUHLvnK3Y/d51q4WRyVd2dHlfujlSXznI3haL8PTvU6BTpcARM19Gyq95e+eu8m3zfXoLc1PNNh08mei63xewF8VSAEZ9dJhZexWbuaCdDaQKmojsBaR8HjkIwagyA4j8rWGI1qK4EfAOf3zJERCn1Ua3omZeYiJfHzrVKpkRqbemHYwKiCwAtgnYv6cFV5dri19YXa497ZY/a7+Qt6/f41Ku8t66xA7Ry6/SWQYXiOiv4QDw4ewXuIjXp2XhRCZe8L4/oPh2P7O3/nv/2Zb0Hom5QKAVGTbLJwTmzUmgVzmh0JTe8THTZVvGBimxpNu6UZ62GazX5mxUfDdJYIyb2VZcIsE4l20qwiFcKYDEIBwrHH4KEiFTkpOgORjRNcnLfxIc5PeAFqF1A7D+sc6rrCuHIoqyqxdSpoBopMYc/qCi4+chCF0VCBICHSzBlxQC62siS9mjB9VbR47pITmk8Zg34GgELUi0uvgQLibI0EKNJYzjMYAXq5wWA4xmA8ghVBYELg+CFl1siNQpYpFNogMwa9PEM3y8AAfF1DK4IxCrYWZIXBeDyCkyj3o8BAJeDACF5gdNSNU4HRyzPwuoFRGQaDLUA8rBVYRhR51AzrHThXEFgMywqsMnS6ObqesHdtHdXjZ1C6ELNaFfUAHQSk1WpV10/rifw5gI0WbhbHL3/wI/5vvOS7Pqu0/5AO2eGy0pc110wIAQQPHUK6FuL1EEFo6lMsIlAce7UOWPEiVzLc5fgq1Mz/9qu/m1GPbsyKpRdmJjuYqWjbbUwOVhqKdXJZjhRqsTXqOmYuzvoNBL6HdTYhI/z0W25ZPrB/z99ysDdlDGNYISu6MKYA2MSSuQic96hqh6oKGFcWm8MBNoeD4Kryfufk94V4klH/X6994eVdg5dyll/eKQqYLIPOI1CHRgszeMBbBOfga4t6OMZwOMZgND4dNocfHYzdb/+t//yhB54s18FTgZjQFIlmyldTUzuROGVPkuT5hUEqFe+Yk6+Hws7OyMKU6xzaa0lMc5ZcoA2INUCE2vvJQKcXQBTBCcFJ9BOhUKOqagxHJYajMQbDEUZlNZEIqa1DZS1KW6OuLWobs50QHHq5Qa4IB/eto1Nk2Le2gm5mgBASsSGVPEKY0LiBGXLFeXTl5m/TnzXqBdKQIARRXoI9jCZQodBLQ6DWLsXn1jrZMESzda2ATOnYE0pK2oqitA6ptDMOBCcAPMGrHKKSzUNgsImZZ1VWECgM6wqD8Rg+IGZ9eQ/kEb1fhha5DSjyHFmWwRPBVnXMTjsGVV3DBYEyGaxz8QWFWNNnNlAB8ACYuA/CdQih24LQefpCVX385Gn3G0u+Pmq6+ZIOtE+8wFsH8QFZ4aFVHA7VGnNs0OCivJb3Ie0MPQKFfYblWT/76ud96m///sdGT2wxDIe7PfOG/sryVd0iQ7dTQBmdbBV0nA9LS0E9HqOuSpTjMcZljeD8Q9XI/unPvf+TZyfH03Qsz9XVmckv7RQ5OlkGneVgk08+XyKNUrbDaFxic2uA0bhGNS4fs+PqEzbg1n/ykURGeN13H96z2vmR1f17X5Qbk2uloEyGLM9RBwsNHbfK3kKcA9kablxjVJYYDofD0dmtT/lx/f/VNtzxZLoGnhoCpiKT1oQ0wphNXpNYYUEi4TaIjzvoiQNnAAUPcNzRC6L9AyT2TqZlqjBn4CCyXama08IcS1NKZXCkUFoH6zyIFergMK4dhlWNjdEYZ7a2sLE5RDkexZ1XiEObIcS+vZcIWDEl4zjIGaLeWSAGKwWlM4zqMWpx6A1GGI4qLHdrFEpFnx7nQdSAT7QTjrYImAGesDMDStkT0PSA5gFoUrILQBQlkImyQwgWxASlAevKyEzs6CRd31DPk/05ORAslHcT1Wqi6DpJxsCHgDoA+coyTp7ZwKjyOLlxBo889CiG4xG0Mjjx2AncedfdKGsX2X4ggNWEGh9baD6WExt2YiN6EYCjh/bi0KGDyEyGLMvR6a3g4JEj2Kws7LgG+3gNsQA6CLTmXAgXM8IS2nmhc8avfvQT8mPf8cx7xNW/rgeDo3apfp7zVdGrOnDOoagLGJNBZwaZKeKGkFVUKrA16kQO8LYGgkft3HpZj64n4f3A/JzOueL/fN1LTY7Rzfly/7tMkR00mqC1BpGKdHGTg5VCcNHE0tkKdV2iqkrYqj6L2t1qrf1oc7yfffMrLj6wb+VvkeZLmQKsc1haXokkoES+keDiZ7quYKsKdRWBbWs83BxubP7peOj+1T/9szsfAYAff9ULltdWOt/XX1l6FVR2sVEGvd4SAiuE4NHrdlGn7EesQ6hrSFliXFbYGo4w2Ni8K4zt741q97Gf+G8fdi0IffPrcQEiYbbctiNLkSk9OGqIecB7IAlsiigwYaacdz7l6unvo57cdA4lcKRQ1lWNwbDE2cEAZ86exWBcYnMwxKCsUDuBDYCVkHTMGjUDQuMtKsJJ2DPOzEQiQ/S3lzScKsGjW3RQKEKn24NSJumsOSiJgDWhnCdxV5kRSp0a9M0QE7a9d3IOdlxjICciIB0Vs4NENiCAqL+FeJ4R4CJJA4h2D8qo9FoYWiuAFMbOYzQeoawsHn38JB49cQpl5fDhT/wZvABZ3oE2GUyRwdoaRIQz1iHulxnOR4Xi1JLDnJs6Gu2/+EIVA/c8ehL3PHISRaZQVx7aaFx93XUgY0DWxYPEFwEKASzKCGQPid/Twsz541984tbxf3/z028z4+p3x84e81i6wlsL76MwbZblyPMMPvNQxkBrg9pFxqLzcUbHuRoED6XN0sqetUs3H9+8+ImAkFJ0uNPJ35x3O5f28gyFMbF8G38LQST0SCLzWFujTjberhw9akv7wZ/5wJ8/CAA//fqXdfasL70jL4qbgHB4qdfH8vI6rAuAzgBlIK6G9xautnBliWo4wHiwgY2NMzj56GNfscP6/4Xq3NacX7ejn91f6b+eO8UNmYllQkpWLlmWo7YVBHHDLM7BVjXqcYXN4RAbGxuPueH4fWUt7/mJP/zImSfb3/8pY8AVJEhInjZCMpnpmS0pBYQon8GJDjpDYNhOppsKwkUJd0qzQD6EiWRPdN2kqNIcKEnWECpnMXYWJzc28fiZDWyNxtgajFC5qMBrfYCX6D0EMgAELvipJ0/jI0SYWhc0bp+J/c1TxIRAkOcZVlaWwUwoihwIieWnpoxsSfV3gUcjeAoAOsl077R+CDu9hmTqXIog8D6CmOLYY2l+35RCFXMkSSBOxRM0rLXIcwOwgZCGV4TReAxfWWyONnFmcwtf+OKXEZRCFQRZ1sGpsxsoYbA1HiOzFYLUMLmCUCxJWhBcmFp3EBOCl0nptSHtT7ztCNAZwVlgZKOM02DgAQEMHO5+6CG4QCitQydfisw8BoL14MDwIn2SsO/6gxdlXzj+YN1CzbnjX376syd/9OnX/FHP4embG1vLRZ7tD8MhBEiUeQdfu6gyMOkNOfjgotIJE4INYAVNyuxVWh14Qguhkms7q6s3dbq9FZ0psGEQAyYzkCRMLBIi7b+KmyM/tPDOOTse3lVX7lMTMkLGl+QFXhQYl/eMRp5lqKyHyjsQpeEkmibCO8BVcNUIoRqjHGzBjkcnUdYfCKJu/Zef/IIHgL/7mudfstw3b1GGn9ZhpYzOQFkOkILWGs7XUZkEgKstbFXBu0j0Obs1cL6ubi9r+7s/8Yd/9siT8W//VACh6KNA1KyLM72hJqFJumNNGWrSaE8Lb5rZCVH+LC3wtLAvMmu3ECjZUEfCNUhlqHzAqa0hTpzZwmNnz+LMxhDDukZZ21QXUmkQlRFEwSfVAKUUoMJkeHWSjTCS2kMqBxKDECDBQzMjzxVWeh2s9btY7vXQKTKwEILEmSEf9SEmGZ4scD9drDcnFyTdkzYA8D4kVlP6o0hToowZHYhTf0yDQHBKYVzVcMFjYzjGiVOnsDnYArIMZzYG+PCnP4PaB+zZdwBZUaCyNerEyCsri35/CWtrS2AlyIyGUhraZKlyqYDQLCoaEBczIiR2nQvwIqidh/MBOtN49PjD2NwcAwqoHPDgo6eRFxrKZAg0gmYDBQJpBYFAGVX4EPYGEQ2gBaELCAu6bzio/s3yen745JmzL8jzbFlrDVvX8Nai2+3CWotADJNlaWaOIRwmBo8MwBLWvfhLfvpVzyv+zh98rDzf8/7UW199TKv69SrPLzFKQXEiIylOiu9TseC6jgs8QCiKDkw+tob4dMU0BoB3v/FlR7sFv8no7PI8N5044pEBOk8ahQwRP53ZsxVcNUY1HqG2pYTR8Mtw+P1/+emvnAKA//2W5+v19aXXr+9f+25tsvXcGGRFEUuEWse5RgpR7LW28LVFlRTnz24OUNnqUUX6U8L680/Wv/tTgR3HRJSnFW+6eM7gCMm0x0ELBDzj0KcAEgdJORCYQ6RrC0130EITNQNJw6BRUZtAJsegsjhxagMPHT+BRzbOYDC2KF2AkyigKkiKCynLYFJRS0o8grOTFEJkOoukJiqpASwBTATFMXtZ7vWwurKMPUs9rPS6WF9bQb9TRCqznxrLTXhwHFlJkQ047XOJbC89zhMWpiVM2Tm4SkBQkbAjnMRwJncVeA9kRQGQwrAqYYoMQ28xHm/g1JkBtoYWZzZG+PDHP4qytrjiumugswxmaRXDzU3c/+gJrCx3kRuDpV4HK70eekUXx44exaXHLsLFlxxGkRt0ig663T601tBaw7CGhGgZ4b1DcLGxE5K8fVlbjJ1HYIPKVvj9P/gv+Mrd9wFa4CE4vVGiqh2kdqDaor/UR0dn8N7DWQ8S32HwPh1BqI0LiH/72Tuqdz39mtvHW/Z3fFEdsoKn662BygiwWQbnHPI8gym6kebDOs6PJWWQCBwKZLI10+09p7TlMQBfPtdz/oO3vm5luadfaforrzCKlzKjYbIcRmdQrLbNyEmU7QkGdc1gY6C00dqYHKiXfu71L7l2Zc/SD/X7nZfobufyfqdAUXQjq08ZuEBJedtCnIWrqmilMBphMByhGo0fHm8NP+yEb2/Or9MtLtp/cP8bWeOywhjkRQcm74CzPDEyI4+VfAA7D3EeTkKsrpSjTeXcx8aV/89/7w8+soMg86s/9BajNfU6eV5ozXDeex+w9Zf++b8vWxD6er9GwooAWmZ27EwNGMkcsRpp1qbRPmNQpFKnjEZkpxW3TAQ6p70VSOwBBQgcGNZ6PHT8JO57+FE8duY0hpWHMEeJeuIIIiRQkhQDJMoyqMaem2IaluxLAACGCUrR1I6a80hpNhr9TobV5VWsraxgeamLXpGjyAwMxzIAiY+JVyq7SfJQir2YMLE/382J9Vz9sLksKBFBqDGLa/paydvJGIPax6zRQePU2U08dPwxPPb4CfzRn/wZbrjxGdiz5wCgOzhzdgu33/4FQDGENXrdPp71zMtx3dXX4vJLL8NFRw+hV3RAPiDTGRAsqnIICgHOWvjgYesR7MhHOriPw7vB2wmwhxDgrEOwHnACYYVMMV53yysABs4OtjCqLX77vf8Nj29swsPCC7C1uYXQ6UaAyxkMzuzI7s1CaEHoCcSvffbOwQ/ccNUfdkiukTzsP725dWQ50+mi98iyVWRKT1S2heJgdEDsh2ooOJFud231Kledec5PveoF9/3dP/jIwkz0773xFjbwz+kvrf4gcnVZoQFtDLTJIiOyKXsnfUkRIPg4eK11Bq0VDma5WV9afs4j9z/4Q2sHjtzEho8Vnc5lhgRZFjOWwByPJQDIgyRej2VdYVCOsTkcYzgcbtrB6JO107/9q7d95TQA/J1Xv7CzutR9dZZlhzMVsk4WmXCU6dhfTdpw5AFxPnoPbQ2wOa5wZmPL1lX5OZTuPVUddkjz/MqPvOXIFVdd8RPLS0uXaoDyIhMPX422hnf++l9557+urL/rR/7Fb9gWhL4eeVCQTJSsE8QImkl+H31jMFXE3i4wSpMMKcniSEjCmKmZL0nmpnFmnVBHI8OroTl7L6i8w/GNTdz3yHE88vhJ1CGqNgchcCAoCDQTcmPQzQsYHWvewUdRVdaMzJhpmS/ETEkzQTEhL3J0iwKdIkduDPJMo1fk6HY6yDKTZnMozlN4DxIX+2EhDZCm8l/si8W5IAJBzxmVYzEZQ6aZpDRpZRwKAiiSOgLiMGyja0eskuaaQuUDai84Oxjg5NlNvP8jH0Z/bR3X33A99h7Zj89+8Yso8vsQxOHooQO4+aab8R3PfTaWl5ehKRIbljpdhOAAcag3zyD4AMcM5yyUir2DuqqSHJCPkjwURVLFSyxlBJ+yIj8B4TxTqKoKo1EZmYDMYGvRIY3veeVLsVVV+NDH/gwPHX8cmgjWWljv0O2tYTjYyjIJa6HNhJ5w/PrnvvzgO59+5XtMWT2NlN5vNRmREAVsQQjBg0PURRMKcXBUAGYDkIcBQFofNt3iDbpynwXw2cX1v/IKz/ovszbPMBTQyw1Ulk/04VSyiI/HD5HZmlTzdZZBnENuFKSLI8tHj/6lor9SiHO9IsvixtDk4CwDiYol/CAI1sJbC1tXGI3GGAxKbAxLjAbDu4ZD95sW/DkA+Jsv/g6zutR7zd69e76/tv7SpW4PWZ6BTJSwmtopJ6q6tRiXY4zKEU5tbmI4Gp5EVX/AVuEDP/tHfzZHVf+VH37LsaMXHfmp0vsbg/c32LKijgicOI/gb9x3ZN8NMnYf/tf/wzv+zQ//6r9/uAWhrxWERAqB7AXihSyzRm80t5YmfbiFB5lffxtRz+2N+ij6Nhl6ZQC1ddgYlXjk5FmcOLuJ0nmYNCegABR5jl7ewZED+1HkjF5RoMijWi9T2kEhzjERRa27kCjRDIZS8byVYhijoQAoIuRaQxsFeJl4J7FHdAsFEghKVAVPpOswaZY1LDg/adlvt4eYfS8aUoYsEDpVicoemrIeMURplM5hOBpjWNZ45PGT+MStt+GmZz0bxfI6vnLvA3jg4ccwGo/xrGfehCuvuBKHD+7HyvJSLKsVBYo8RzkaIiMFNzgLZ11ULwgBQaLymA+RlBAd5yRJI0XWY5wjCphQzL1Pje4QZY0g8CGa2hmyABOcraFdrL/3lIIogxd/5wvwpXvuwac/93lUlYXKNLY2BjBGKUFY8T6YFlaeeATWXwxl/fFs2dwgQoddsGBmOGsTWzUyVqOsFQEqbnCYk4qG0ntW96zfEEr36p977Xc/8H/8lw+enT3+T7/5lgMZhx8sVlZekLF0OoaRa4XQEH8aMk7aZLFMC9EEBU0ZAgsUGJJTfrC3lFsboLIAozj6k6kMoAyg6BgMCYCzCC7OF22OhtgYldgajs+Wg+qTlac//ZVPfakEgE4nP7a+vvSjppPdlButmRRYRz8jZoJQQEilee8cvLVwzqKqLba2BmU9HNyKGu/9uT/51Jz77D995+sPra8v/w9e8XO6ve7VSjw6/QKZ0RAPFYy56KzgYFltHu4WefVP3vnG//uv/rvf2WpB6GsCIb8qoIMgypqu/mTCf2ZzPx3QxK69jQlaeYHwdk8eROq0RFkPJoYIo6oczm5u4dTGWYxsnHXRykArRr/bw+F9B7BnZRmrS13kCsg0wWiGMgylVVRUCEhSIQk4aErhIop2Dpx2bUjSOYxoaCWMdLF6NII/swqsRLzN2nvq5BqQWDyzFuKzoDsL0tNHzwFSJJMznPfwyavHQXD89Bncdd+DeOz0GVx93Q0YWo+PfvJTOHV2A6vLazh26aU4duQwLj92CPvW15AZjW6Rg4KgGm8h1CVQlfBKoarHYFaRBeddskf20z5VWkwCx/cheD+xiJg97wmLJbqAwbkxIA5GA+PRGBIIvbyLM1tjMDSMB4puHxcdOITRcIwv3X1vnNFyDirrqhDqfghtJvTVxL//zB1n33XTVR8K1r4sGHXIByHnHJDl0+uw+aIYmlTcRBFBJRap6ncPd9dXXlWfOP0pAH88e/ylbnZDf3nppaz4QEcROkolLy5utqORhDSxVUmbKtZA8OCGQEQBGQiUtOwyimU8VhlseqhihnM1DAHiK0hdoyzHGA0rDMra1aW703v1AVZ8AgB+/Jbn08pS8bo805fA2W6n10NWFGBtYjbI8dMZnKQepI0Z+7jEoBzBl+UDYVT+R6Fsbij1H3//a/asry597/Lq6iud1lcbBOSZARRg6zGKKA2ODikzgr6YMvUSDu4DAG5tQeirjMv2XaLKcnhImA8RwBwCSElirSUDumZxFU421LODlmHSvI5ZjprotU1mZJCmCEI0cCMdl/qofkAYVh5nt0oMB2P42iIzGsu9LlZ7Pezbs4aLDh7A2lI/KnWLSwsg0HCtiQikEXtFSdcusEonP5UuCUlMtNGkgo+2w8QxMwpQEHEIiZAQ1QcErHXMUnwAM8FTw8ALAPPEpqGRHwphpyGeMEF8SEA9BfNYhov390JwIFghnN4c4b5HHseX7n0IG1tbWN53BINRheAHWF9ewXXXXo2bb74Rlxy9CBk72NEIwZbYGm5BKw0EwelyE0qb6LrpLYgVynKM2juwVvAuzh2pZFkOkWSHEYUeNUc5fkZUpJgAkggk0eE1A94LbG1R5AWc9RgNB+hmOcZ1QMEKIhb7V5aAyy7DXXffDescCAbOC0NQBBHVQspXFw7qC1xWHwm94lofsCd4D6XjQLZKNu+GkwOYUlBaRzt2yuBcAET3l/etXWG0+pF/8uaXjUTk03/tPX9S/vJbX3ak11HfR5qOGSawIngI1A5dyOm8GMiDoRHgI9eVAGgTy+JK4Jwg0wokKm1v0+cy+ORxFUu83llUrsa49hjVHta6BynQHwXiD//yxz8tANDr5jd2C/MCY/JjnSyLQ+cmi6QLZjBSqd5Gr6Da1RjVJUZVjcFgcEr78Kcg9bF3f/DTE5O/X/zeV+1d6mZvKJb776yIb+xojsO4EJAXZHkG9oCzFhws+plerpw6lrNc2YLQ1xa9LDdPH0lYi+l11DTzFKLtLSfiQRJD9GnBkmaRDgHBO4CypCSQlliOO/okH5oEAwMUZYA4gA08MbZGJU6cHeHEqQ2UwxK9IsP+9TVceuwiHD10EP3CwJAgYwedbH2NzpPcDcWUvuk1pRKw0iqeb2zpxF5FiMQEaTIh4UQACGAVFbwDHCBq0tti6NgzCY0FeXw/ggugTKMOHkbFnhYn9l3DaANR6uvwJAkS5kQR5MS4k0kVs+mnVEK4+8HjOLk5wj0PP46RDTBZFx/+wMeQFTne/NpbcM3VV6DTMXDeYXz2OCpbAz6kGSxg5KIahPWCcb0FC4H1LtqC1zVs8FH9gmK5U4UAzQoqU0kglqMeoABKCEZpaCCKoTJFk7y0vbBeIEFBMSO4KLGSaQPrHTRF58+6cmBSWFvKsbbcxebYYnNUQsDsfMiFQwtCX20wnfTQtyHglIXfAyLU1kHnAaIiKUdpDcOxLMVRkj7SlpVEPoHwYV7tv2Btubty8sGH/+yXX/fsrywV+G5T6BdRrg5qxUCmETgCGafPNQLg48BdKoVHcg1L0oH0klijqWynIvQoMpOsWjFin9LGHpZzDtY6jMY29YJGQzcsP+Rt+Lf/+COffhQAfur1L/mOQwf2/r3e8tIztdadvOgg6xSgTEXNIKUhPgDWQioLV5cYjrawMRpiazyqy8HoM3bsfu0ffvD2iejpP3zLK7O9e1d+dHml/3bPuC43TDo38ExQYCgSuNrHz5WL7sNUVyBb98i7PT/3mhcZALYFoa+mrux9YcVdLJq7mHFTRerZzJDQIDxTckNIGQRPvDYjeyqASKWKVwKu9BilknoBxaFUGwSnNgY4tbWF2jl0MoUrLr0Ix44cxfrKEnLDYKmjz5APcEJQRsF5B5VlkeqtTPIJIjBFeY5a/OS8rXXwPipmR222gOBDPG9W8CEgVH6iEkFC6Pf7CM7DSbQXrm0NQKC1gQtRRYCChwZPVLbhKdXIeZLohEbvSKLcT4CNGl4zdNn4fit4D9QCPH52A5//0l1Y3X8Qp85u4r77HsDhffvxule+DNdccTFWlvqoyxGG1RZ8cNDMsOMxgvMQYgQwfABK5zEsa2wMx9gYjlA7i3FVw3oH52OtXCuGZgL5AMWELM+Q5RpKRwJIJy/Qy3LkykMDMARkCjA6ETiIko0AQGiEWRslZ56wnDJtYOuoL/eMG2/E+z/y0ZRFe0jwTPDSoslXF79x6xfD259x5Zfr0fB+7nau8j4ghBlX4mT7rVVkirFKmXyQmDHVDpoVrOAovO3vufTotb3RmiVWfWTZviASN3U62sUrFaWjaGaWMIQokJp0NFLxIVZT0DBXgWTiOFO6a9YXxJkgCemrCGpbY1yVKM9u3m8Cv4/BDwLAP/ieF+87eGj1b2Yd87QA2p8XOYpeDyYv4BWlioUHWQexEYCqcoTxaIThaIjB1tbxYOWDztPtczvxfu95psheYZmvKIxWWiXFFUriwj6qQZSugq9KsLUYDkeoR0NfjsfeOvcNvYa/rUHI+5B5hD0inDHTtOE+I7bZ1OSo0WxpGFwUMx5OhnAEn4psUTom5kA6lt4oOYMSg9kgKI1x7fDYmVPYGo2QdzJccngfLju8H8v9HIUS6MbJNJX38m4Raco2wINhQ8DWxlkQK4yrCmVM3VFWFcAUFQicg0dImmZZmiKP8y5MnBrzglFVAUQYD4bodXvIM41MMzp5juVeF1oRtLXQDHSKAq4qI9khTecGNlG2iDkRAqeGFqEhKyRZo8QPjI5IIhBSGEvAqc0tPPDIozhw6CA+edtnceKxk3jaddfgphtuwDWXXwYtAZtnzkT5efGwLp5zNS5T9sqofcBwXEZK66jC1riMdhUS38NoQwEE71E15xkk2kSXNYRiybHQGkWRo5/nUZXbFOhmCkYBmiVmRUk9vSmJNr2uSFvHZJI/AlWk9R/afwAihG6nQFWVUN4RQ1qL769pJ4njdljeaYx5rguy1OgUNuMDSikYrQAmsFFRHCuV0MYugJWCyQh1jVU22Wqv248bN1tDISR9OErkGoCbv+/2oWuZt3GZ7Y/STHcxqppgMlSOtIF1LpZ4q7rGeDQGeW9NVd/qvfrEP/zopy0A9Jc7N/dWeldAmaPdokDR7YK1gU87v6hlGHuOrq5QjUcYDTcx2trCcHNzKGP7iaq0v/kPP/iZCZHg3d/3uiPr+9f+J1MU12eaO1mmJ5UUCVF524Y4NyjeYzwaoRoNcWZjK7jh8OTmoHz4/3zfJ9zfbUHoq7x+g5jA0pt4YWN2wHL6vUzsGDgNXgJQM4oJSM6rJNOrK3G4JTXehVRkU3H8WWUtxuUIPlj0e33s37s28cBRsR4G71IjlAnjcQ0X4uDqqBpiVNV46KFHsDUY4Ct334sTpzeieKn36PS6WFlewcrKCvbt24f9+/djpZOh2+kio8hFc9aiLuMivVWOsTUY4O6778WJE4+hrktAPA7s34MXv+iFKFR0Cz24dw3lYIzlogMKDlrFbErSzBPNULW56VchstEUR2HREGLxD0k3zhLh7LjCYxubsBB88lOfxpfvPY4XPv9mPPMZN2Hf6irga9iygtQValfBJr+Y0tbw4Gh25x2G4xInz25gczCOyuE+wAtNRFyF1UTNQik16fExVNqJxuHb0nrossKW0ujlGdb6S/C9LgrDMErghaC9j4OtSjU6SHGQOchE7inPcpTWgVmhkxfYrBwUEbq9Hja2tuAldGhqZdXGV8Uswqar7ZcYYSuILIU0TN4AUbRkV4CK1uyQ6IhLiqF1HGtoFBBCiCrGRIgKGip+VryfSm/tJDYlrzGJWdjUYG+epEOzUiAyzdYifvHEkFIbg06nwObZjUHHqLsq4q1YMnvF4bW9Sz/o2R3qdXtU5DlMnoN0BigdN1jBJXuGGq6sUI5GqEZlFHAdl49Iad9HpO9qzuvnv/e1vQMH9/1Qd3n5BmXUfoMArRWIOK4l1gPc9L8lEhzqGhujEcq6erwajG4f2fDlb/Sf+Nu8JyQMkI7XCM1kHokPJbNu1jOlOkxlOhr/n0AzCj/J1puaEg1P3Ux9AIJzGI9HYPLod3OsrfSxtroMnZmoSpB27o4Yg3GJUVljczDCg488itMbUS9LFTm0Meiv7sHeiwm+cwpbgyG2zpzF2UGJs8MK5uQZPHryDNYePYFOt4BWOr4Kijsya+tYh64DhoMhTp0+i5Nnz4BVwNrqKnzeQa0MHn70IYw2N3HFsYuw0uvi0No6ljsdSDLhEhLMOYojCZOSxEawxN+HSVM/6o0rZTAqLb784IP48t33IsszbI0qHNy3hssvvRh71paQkcAOB/BlCfEezteoagtFGp4JFTzOjqMfytZwhI2tIcaVi2VPxHkJSTs7L5FIwKm3BWIIq2i3AICVgWKCdRY+CJwEWF/BB4L1Acu9AkvdPMoGeQcdLDIjUBTVlKNnTSzNMQCXxF+D93C2BkPjmqsuR+UIG5sbCIC5QM/DNnbFIKmC0P0Ab0WFeJpc44kMF2najGj4KGrSvzQmi8PHzkWDSk3wwUMpD0mahs45cLpWmXmOWDOrCNIY2TUZ2KK57anE1wyRR1TctLBO+1cPYzJ0Ox0ZMiqjqPuz3/OSi5dWuq82RXZtVpj9WaaiQyoTSGsQq2gd4lMWZOvkGzbGuKpQleMNquo/r234k5//4G0CAD/9+leqpeXui7or/VdTbq405JHpKP4KaHgPWBE45+LG0dUohwNYazGqqmE9Gn1qNKx/15G6twWhr+UCFhGR4AGRSJumOQXoubEWCXMDqzIxwElSPkLwQolNFfsjFOLFyCEaeGdaI4BQeYd6NMJyp4P+8irW9+5Fd3kVgRhBgIdPnMSDjzyKja0xxnUFYUJWdPDY4ydx/4PHsTkYIOtkOHD4CPbsraFIodNfxmBcYew8NjcHsCHAAZATJ3FsdQUHDuyDcxYCQl4UyIsslRWAYB0oePR7HZw49ThqF0nc47LGn996G44ffwSnTjwO1hk4eHymdNi3uopn3/xMrC53wCihIFNbh0Q0iE4YscQVN1ORFBBdVKOEyv0P3YfPf+kuWC84cWYD+w/uwXc862ZcdPgIfBlnJTgJVIq3CAGw1mLsKlCW42xl8fjGBs5sbGFYVbDWR7+lVCb1IrGhnIaPjTHIMgOtdRSMFYLzHmVZJrfctBARIydEN8vRGFVdw7oeBMBSNwcLwXNAkBqaw6Rf0Fwiihi1t9DaIHiBY0Iny3DowEE8duos8jxHXY7ZC1piwtcQ/+Fzd/nvv+rwGQTZ8j4kS6rGWj6Wy1mpyHxsysUMuLoCc1RVoLRBbEwYIzikjEiruNlkhvcBxDpl9dvGEcK2WUHsnJmj1Ef0E72VVE0RlYSHAaUEnU4Hy+trK+Ozp28hG6xZ6uxZP7Tve7zC5XmuUeQFjOmCdRGZuCGqvsPX0b6irjAcjzAYj7A5GtaDsxufDWV4T4C5NwLQK9Ta2tILDxza/ze94hsMBe50u7HErg0YBs4GiHOovUVdl6jrMcrREMNxGcYbZ+/cenzzPznJPvruP/1E3YLQ1xAEWAKNJQQvRKbxj4linzTxk5GGeJDSneb7qU9O2nU3VtUhajYhZQIaDISQGphAR2XoZQVWl9fR6XfgWOOBx07hvgcfgXUBp8+exiPHH8PGZoWt4RaKIsOll18OnXewtGcdm2WF4ye38MDJOwHciYPrKzi4bz/WVpZxaN8++BDZfYUx8Kxw/VVX4pJLLoJ1FooZeZ5DGZUsE4DxYAvVKNpE3P752zGqgeFohNLGobm9e/bi+PHHce/Dj6HcGuD0qdPYu7qOE5slXvyi5+LwWgceNQCd5nETW4h40phFEiIlHTNEbx28B7587wPYHFa46VnPwp9/8uO49NgluOKSy7F15iR8OUSIvRMEH5lD1jrorIAnYDwe4/GzAzy+OcTWcAwXEgClRQUkyLIc6v/P3p8HWXbd953g52z3viXX2hegsAPEQhIkJVOiTGqXZUuyZVlqu92emA73dEf3dEfMRM90xISnJ8J2d8hjS+3xeHpshVpye9TeJFmyVi8SSXERNwDcAYIEQVQVgNor17fc5Wzzxzn3vpdVBZKyJZsE8kYkCpWVlfXynXvP7/y+v+9iDCImzURRGIbjEmMM3kd0MeDI0aMQA9ZZBDCZTLlx8yZ1U6OVTl2Rd/gwIxAJcY1RqZEydUTOB4r8ACdmVNrMlFK0ziVNihC44Jns71PPZ8QYcaBbF8rDUvLveJgUcu59mLaZoRhckk2ITouW9S1CqcymjhSm7OeVg0GRRJ3eIUKCVGMXXJkPFsvzvjtBcogOis1Q7526IEhC1xCW4P4FhC2y8WqMMBoO1H1vfuI9Rqq3tt7RRNZWSqNHQ0NhCrQZIKTB5llSchFvaOdz5tMpk3nFflUzr+qL3vJbNsj3//SHPpko3ivDR0+cPvbfovUTQ1OsDAqTfgadiReIBDPHgLMB1zbU8xlVVTHfn151+9Xv+iB/96c+9NT+v4/1fX3DcUJYQdyD6DqLhNgp/Dtngy6qOxuRijxW7zz9RexC2xaMM5Xp3lIEtEjzBqkUISSIRheG8cYm88bx6rUtrm3v89Llq1x49Sr7kylra2NOnDzNibUN2lc917b2ufrJz7O5Pub40aPcd889PGIMPkY2N9Z47NFHeOShBzl+9Cjj0ZC2avAuMCyTV1xVV7RNk2nMLgnZYsT7pHMar42RKyPi6WM8/MDdDMcrTKYTplWFUAahNL/0y7/K3mTKpKpxQrJ55iwf+9znEUbwHW97hJPH1lgdl70zhMhD+w568D5gQ2ILSq0IwjOd1dRRsj+v+eKXvszuzj7BJ8JFM52CrfFtRWubRIOO0BJoraMNkb15w829CTvTCucCPvrUjUiRaNdaUwxKjE6stw5aCd5SuxofYMVoTh0/ykMPPcCRI0cpyoKdnT0+/9xzPPvsF9je3k6QRIR56xB7s+R6LIZomQxivXM4keKlY1gIF7XW+Hzuba1DFAZjNOtra3DpMiC8D6wclpF/1+dYzUBNA0QfkldA7DweY2fZk5/phMohjQGfhMkL+kCKfNCmQHiXoGNiDmckE1HkHckHkY4JKg5kbB0oQCKlpHbC9+6/izFA+nOlJMPhkBCDaprmiDYaLSXj0QitTbK0ihIfXNYDtbh6TlvNaZqaWV2zO5swq+pLvnG/Yb38xZ/+0Kd2AH7qx3/w1NGjq/+1LIonpeDYuDQorQlS4mMaRhspCd6jBSjhEDEhEfPZfOonk6eqWfvrf+v3P/vvLYzxdV2EpBRWRHENaDsxp6DbQBdzoGSoubhVQ8i2Oz0ryhNiyoPP/XXSE8hI29aYsiQqiZcC6yX7s4orW7tcvrHN5ctXuXRjCzEcsnHiBK2A7emMJlxhPBwhteaBe88xKAoefdODPP7Yo5w6cRyj05C9NAVaSxSRWE+YVft4m4apLZHoHc7abGMSEyMu+qzPSfHHMrs4xHyKq/d2CECpEt6sROQv/cSPsT2Z8MnPfI6PP/UML196hdH6Gp954Yu4Zo93PPlmHn5wBa0UhVI01tM2Fc55WuuYzGZUjcVHgTIluijYnc4IusQUA15+5VWi94wGg2Q53zREVxNtg/ctMSosIIsBrZdUbcP13V32p/MUBpbnaOVwSNO0KdzMmERbtx5pIQRLYVTvrWe0YT7d5aUXn2dUKlaGA04cO8qbHn6Yhx5+iHPn7uHTn/4MN25u0czm1NN9KmvZncwhBMbFCsWgpKVNdj7eZcquTDY/wWdtSNqYBmXSXq1vrFMUBaCUUPrUW8/caz776gV7WE3+bedCYuZ8mJdCeuusDhk+98Elz78YchBh7pClJMQkMFdC93PdNJBPMgIhZD8bzgYZPXHltUx7u3nQskHvrbBd31HJ5GASQk7pjcl/MoTkdxg9ECJlUaTCqHW2Sy7SjEvIFPQYPMG1uKZKyattw7yp2Z/P9pvZ/F/6hp/96Q986iLAT/7Z7x9ubI5/Yrw6/nalxF1pvhlTQUNhTNn7Jqak5kTzTjC4t7Gef3G2O/kXUahP/ftc39c3HCeo8fEiIc5R4khixsiDgJ3oaQrZwDOiQkDqpWA48qlL+oX4UihcBFkYvFa03lO7wF7luLK1y9OffpbB6hrzxjN1gWZ3woq1ONsyHBY8dP+9PHD/AygReej++xkPS1ZXxqyNVihLlW8+TwwNsYm0zuKsxXlLcEnzIwDn2hwTnCEKuuyjlEwpsrDTuWTTI0WOfyDl6khT4KTGjEasForHH7qfjfUVrt3c4aMf+zhHjm7wwiuX0cMRenWT+8+do7ENN65tsbu9xXQ64+VLV3n18lVW11aoraexns2jx0ElrdPxEyfY39vlzMlTbKyu4ZsW3zZE3yJD0l+5CKoYErWhrht2ZxW7kxmN9bgQiUEyGI84d+4ednd3EUaxt7tH26aMougdMVoYjXoGlNaKQgtmk11efeUCInqMhLNnTnP65Em+4zvexYMPPcSFl1/h+c9/ni899yyzvT2quqEQ4DdGFMagpaSuG6IPKJl09T7G3vonQFKcK4WzFmOKDNl4LYVcL9Pg4bAI/VtePkQ3mUxn5crYe++1dw7vHEGnULuYBcp5SJk6mhytEmMgJJvepaIhs/h0WRMU+0yif9dNZzl/WGYCd8h3Sx6lJr/GPLSVnat8fs0EQZCJMu1tg21T7Ld1jslsyu50hnfhxWj5pz/9e5/q2Wsra6O3bBxZ/VFVlg8Oy6Sf8iSoUimdJBY5rTYER1NXzOcz6rbGVrNronEfaqP40P/zw59qD4vQH9oJispbfyHKOJFa9bPFTKTp54y98aYIPSCnZEotTI4FIETyXovBI7TGE1KUtDHsto7t/TmXt3d58eWrCDPk6t4MP6nToL1tsK3nXd/6NpSM3HX2LPffcw/Hjm5SSEmpFOVAE50n2grbtFjbEpzLzgcKT0y6oOCTej+k1xxCcoUOIRkk6qz4dj4VrQi4KHGZAahF6nzI2UlSSjAau3uT1fVNxjry2IP38sD959jfucaLF17h+PGTfOmVa+w1TyH0gFcvXuDlCxd47NFHuL435f0f/SR7tWVjKJnVgTbC2uolTp8+zT0PPEDVNNjWcvzYMUpjaKoqebs5m5XuiiAVyhiaKBKlfF7TuIDzAescpig5e9dpfvRHf5TheMT2zg4///M/z3Q6RwgoVOpu51WFrAXGpKH0eDDAO8f2zetUsymlKbj/gYc4euoMx44e5fiJk5w+excroxG72zd5YWebYZFIHdVshl8bMBoMs09XyJ1yhlyy7ghEStQNkVcvX2W0vtnRF5SKYb1EDIH6sJz8210hRl9XdZPsSCijT/d/8CG5B2TbpbTByyX4LTlEhqWupdcDwiK+JNALupc9EQ/AbLd87tYQS3GLm373baTIjo3CJ0f8pS6t0+vILpcsSIJfkKS8a7FtRVNX1HVFVTfMast8Xt1UQTzVonpR6k/9+R8+ceLEkf+iHA8flpJxEvAm2rlUiihVCuOLgRAsITiqqmI6q2jaes/uTz82r+2v/uSHPnPh3/f6vq6L0Cu7l8OxYmObGHdiT6jJqmYpby9Z2a4jxlyE1MJNKg29C3xMNFEXBLIcsF01fOq5L3NjZ8J+43j5yk3KwZh565i0NWePHuFtTzzKw/fdxbe+/Ul827KxNsZoDWGRBd9OA+Rha4oUCLSuJYSIj8mBoXUO75No1bkEQ4S4UPCIDC0oGftBvbMWpE5wogAvPVqkaAUZfarGNp2Wdm9eQxhN3dQMxyN+4LvezTM//ffRg1UG41UqG/jcF15g6/oVnvn409y8sUtZKu675xyl0YxXRwShmVcNX3rxK1y8dBllNLt7+8QYKAqTCAK2QQbfe9RJlezzpTJ4G2kdTOct03liw41WVvieH/hennjiCb73e7+H9SOb3Ly5xYc//GHOn3+Jm1s3sc6jjaFuWpQUeR42hRgZDwd4H9jb2+fq1atcevUSK2ubqLIEFRiPRjzxxOOslIZ/JQTnX3gBEZMuKPjk/TUoDdb6PsBPyORiYRubMHwlcD5w/cYNhqtrrK+tUc3mAz+r3jbf3/3oX3rH4/HRB8+tro6NkILdqm6u7c+qG//Dr33IHZaZr9lexBBjq6QKQsglfz+ftDPBoYJfQjSWDpe9k1vuQGQXT0KvdQsi5lzI+O/cCXVkp65qdd9PdW4LUhCdzFnLMUkYo+j8rfC2BQUIj7OZtVZXzKuaybxmOq93tBO/1zbuF37qfU9vA/zkn/uTxbETR/7jlfWNt3kRzmotEVolKyKRoT2fiRzB0TY1VTVlZ7LP/mxWuf3JU9Xe/J82LnzqP8Tqvu4dfqVSu9676zEGixBF7F0J73jiSkK3ELI+UfaFCQTeRoTS+CjxUjKbNjzz+Rf50sWLzKwnqJLKwc7ejDc/cB/333cP9919N/edOcnpExsYCXVo8dMJdVv1RqPloKSp696Cx0ewzicrGutoXGAyb5g1dfJHsw6f/dm892ilKYoULy0FlEWOhDAGIYs0I4kBScrWQXampFny5ANCC6rZDF2UCGPZnc/YPHaMd77jCZ7+0suc2zzO3efuoZrNuHTpEvfecw/rq6ucOXWEhx56KGUgyRTiZwO8+fGHee8HP8oLX3qRYphEhPOqwjmX4ayAEcmQsShLhCmxQlLVWRM0mWOtZ2VtBV1o3v3ud/HwI29itDJMGiyleMtb3srO7i43t3ZonUUoSYgyaYxiZFa1KK0YlAPKYYHyMJvNufjyy5w8czdHTpzodivWVlZ421vfylph+PRTH2f3+hWK2DIoVZobdFHPmTXpQ2ePlB3MMx1+bW2NVy9dYjReIbbNqIr2++bTG+7uu55YffOTjz44KCQyuMl0b+/S+YuXf/6v/NB3PPOTv/2R6WGh+aoIF1Ion+C1TBTqCpB3eOeROScqLolOF+VEpi4pmxkmBCCxOftgyyAWBATuTDr4Oru2/C/mFx5J3z8mCC6IkLwnvcj+K9ltJXYO7xbvPEJ4WltTN3Nm1ZzJfM7+tG6q6fxTsQ3/sHXh0wB/7Ue+T6+tDn9oZW3440GqR4amEKZMEeVRSoQ0ST7hHIqIbWvm0332JnvszGZUe/svVjd2ftmhPvA/vO+Z6rAI/ZGQE2QlkddCjG0K90gYPiEJLOUdc9pCz34JIYVfF8pgXYpT8AFmleWLL13kc89/BWcMkxp0KXj44Uc4urbGH3vzY9x/12mUbxkPFPXWTWrSBjbQmlKK9ACFwHx/n9Y7rIu0PlC7yHQ+Z29/zrSqaK1n1lhmVU3rbE8yiDmOGwRGqewCHCi0YGU4YH28wmhQMio0hRQ9mSLJHgJeLQS3oW0y3Jh0RTEqqr0Z73jyW3ju4g22bt7kvIS2mmGE5Lvf/S7uvesURgiGpSYETzWvsN4x0IbHzp1i703n2Lp5lcrVlKZgNp/hXEspBVFKjE7xzEUxRA+HNLOarZvb3LyxRdNaTp46hccSZeCjH/swVVNz4vQZQkjU7AsvX2B3b4IP6VaOUYIwhCU/5KrxTKqKwXCctDsucP3GTbZ3d1k9eizPx7LA1VruOXcX0j7JS18s8fMdsFUfCZFO1ll9HyPeupTwqQsCkrmzfPt3fDvv/+DvM59PGRs5xLH+1rc/9qNvfsdb12bzWbm3n97nqppfXtvcOL21tfd3/9vv+db3/u33Pz0/LDevVYRk0FrFgwUidUPBLwIJo/d9hHx/wsodTzfzSZ1RehZCZjpKZEpolbEPsvx6koSXYbjbMJXOYYNuTiv6wLLUjUlCiIQgOkVRml/5Fu9bHBZrG+p6xrSasTebxvm0fZXK/roL4vf/pw89Xf/VH/pevbE2+oFTp478FaWLx42UQ1MUKKPzATwxOpMmyOeuako1mzCdTahm8+vV7u6HG8fv/eQHn9n5D7W+b4AipBoZw1UfY9vdK4luGZLwlEVL0ItVRY8m59ujG2ZqPIpp3XJ5a5fnXryELErmtUWrgqPrmzz52GO85dGHGbiGws0RzRx8tpvP9iFtXTEoB3jrsdbSWEvjPU2QNC6wV9Xc3Nnj5s4+dWPxMaYBvfc51C51ElGI7BYQwHlk53HlA7uTmsmK5cj6GhvDgrFRxFJjhERmBwTnXXo2hMwO4jLFF2cRbts4BuWIlaLg2s4OL+7toETg7Y+9iTMnj1NI0NHhphXOtYjokbbF1+CBIyPF0bWSa3PHeGWUFOo+pNgKmdzAjUnx5hFB4zz70zlVY5FSc8/d93Dx8osgJU899RTbu7s8/pa3IqXGOs/nPv95btzYToalWmN9QAmdsPXo0abABU/bOryPRJ1Ws7WO6WyGczaJWmNS1ZcSZnXFdG8HfEOpDc61OcETQqh7OrCMkihDMrOVEqMLbl69xCNvepQPfeRjrI3GbChY0Rtr3/LWN7NqFM4HmpDshkLkzNzF0WB19T+fTK5eBz5+WG5e6xkGJaUSMUrZb/rdDCdk13mfolcQIHW23MqdT1iI0hP7TUF/0ExFID1Zi6TL1ypAy3Og1/rzg2KjTl9E/1oQaU7T2X7hWQRPxpDZag3ONrSupW4b6qreirX9fW/je3/6I5/eBxiNisc3jq78V0LJR0ZGDrXRINJhTKjkGEGUNG2Fty2+SYanjW2oqvk0TCdPR8dvItVL/yHX93VfhISUjQrqUu3aWpmkPpYiRQ50Bh2CpFP1nQ2NdxgFpZIo0Z1aAl5Ai+Di1jafff48k6ahcYJgA+9+1+Pcf/+9nDl2nIGv0LZFx+TAHJwjSIVUCdlzITKbVzTWJ9jNeWrnaBDc3N3nxt6Erd0plbX4qBLzzWcqqkwkg9iZleYHJgSfvLB8YvI5In5WMbeOba05tjFmY32FjWLEsJBE26IzQUHmcW7iqaWTmo0e52qMNrzj8Ud4+nPPcenGTc6cPolD0FhL4RtisMiYUkyj8Im+HiPReTbGKxzb3GDHblMWJdeub7F/tma8uYESDi1zQpIIBBHZqyomVQ1acXT9KGfPnObKtfPpVNi0PP+F5/gf//pfQ+iCumm5ev0azqVdyndDP5lgR3K0hIwRFRRGGKRI6njrbBKUOoeIyUVbCTAxsnvjKluXLxHbmihUfkQs4CkktL5BaUXyG9cgDBZFVbV85rOfZWt3Fzvb58TpI5xZW+FN505zcn0V7V3aHFB4n2ZL9bzakFq9eVCIn/jPnrzv/M9/5vy1w5Jz+6WkUOvjcak1UolFtxJECkh0wSKdRqsSoWV20Ir54JgWV/YEpGyvG/O0SISs/RIL2vYyXJ/JDMuEhP7ceodCJOmcRBY0boTos7akUCzkIkkKErInpRCBmJOPiZIYNU0jqGo7EdY9hXW/KGXxKsDf/HM/+MTRE6v/vRmvfJsqzKo0hqg1aJ0o30SkT2QZo6CtGuo2aYz2plNn5/Pn7Kz5F63nYz/5e8+EwyL0R9vLV651LwXhplKbW1xxPQLVi9yiCBkT9igRKeQiD0eSvP6v7+5z/uoNru3vYduAdZF3vvVBnnzsAU4dP4om4qY7FFqDTzBV1OlGDNETfKS1FmfBBZhay7Ru2JlO2ZrMuLq1QxsjcxsIUfYRDZKIlIrGZT1QDL0eSGbxGVH10JG3gdZ66tZRFZq5tWxP5zx0392UpWY0GiGjRwSH8J4oU3ZQECnWQnry6dDyyH3neOXyZS5tbSGU4eVLl7i5vU0xNCglkSrNSlxKEcoD/cCoHLA6HBJsy3R/QjtpaWxgPF6HKqKFRSqPj4kBd2Nri2lbc+bcPbz18ScZr4zTzMUHRAzMZnM+8fGPIVRJ6yNmMESroodAyBCLlxlmDVk/4nPon0gnZp8NUiUBQ8oSmu7sc+PGNa5eOI+d72MyU1JKA8HhY0ApKIXES0UbI8qUIEtMMUY0Dd///d/Pr/zSr3D3ySOsD1MXeOb4UdYGAwohsSF52/koaBpLqGuqtrkbLd4z29/+8F9+2/2//g8+/dKh4entnZApC6W1jKkIkWPiEenwGBJhR4eADInajMrzmCys7uNYerZazAWIJW2Q7L/m4B5yUDN0p+LTd0d3Wr3lCOc8BWIpyTd1RJleriV4RfAhMWGlgSBv+ln1m8Hr56Um/vUf/u77N48O/8rmiePvRKpjg0GRXEa0RhiV2L/Bg00wpYyOGB21s8xsy2yyf77dn//reRt/+2/83mf2/kOv7+u+CF3avRSPFke2BXH/tra5x+AkvdcTiR4pc7h8iElwZvHMpzO+/JXzXLt+E+sicxf5Cz/8/bzpwbspZCS0Fa3zKCIqApl9FkkZJwkaaplXDS4oWh/YmVXc3N/n1WvXmDUttXOgy96iLQSfEk+9w8VETZUqCeFWV1aQSjKdTJJpY46uCc6nouA9XmnaRlArRT1XDAqDPnuc0fFNCmkQ3qNIf9e5pKgIUiBdKioiBqx3EGNylTYF165dZT6dYMUIXxbJEl5CUDFRZtOQBiEFR1bXWC1KdmY1KM3OdEIrIsZogm1SXIQPtKFld2+PRx5/jHe+67t55P6H+eLzX2A4HDKbWaQQaAmDckgQyeBRSpVneykGPXl3hWwwGpNgUAtkkULt9MCkoq0E5UChRMA1U7a2trh08Tyz7Zu0031Kk/UUtkLE1A0bZVKWjZQEBKowqHIM5QrPfenLfPFLL7A2LJhMK558071sjAoUie00HJiUQZMp9nVVM9ndY2f7JgGkDf4+NRDvCYSPADcOy84d9nByxpNMrged3q8jKoTOjifEPPyXCBEQyBTt0HUuMbJsUnpr4bi147lTsfl65kLdn936ffp9hyXaeGdDJVO8gjEFypRIY4m6wNeN3Hv5lYnWhuHQ3Ld5ZPxfrx4/9h16OLy7kIpCa7TWKK1QWiF8JOKIApyzzJuKuqmp2prZdHrDzpr3TWbul/7WBz9/9RthffUb4SaWSu/K4K7EGBsQZXdrd0mhnU4o5tMQmckihep1IVIbrA1Mq4rtvQofwQB3nz3NuChp6ymtaylEmg/EmGIGpE4FzjlP0zbMakdjA21wTBrLlZtbXNvZZmYttXWg8oDSeSDZAq2OxwgpqOsqQ3CJraVlsgEZliWxSB2B9x4vHUVR0LYtdV0DChc8Veu4ev06RkWMlmyMh2wMy+yCneAAhEAoidWe1lm8ENTeJVdpqZAy4dq2bmgGCkNgOBxitKYY6ITLe4+3nlC1nDlxktNXttjdfwVKwXNf+RKnzxzl3iMbEFUe+AdcG/DW885v+w7e9e53o4Xh0tVrbG4ew1oLwhNQaOVwIaKlQGuDd9m9QkSUkIgMLIqQTrpCaQbjkuGoYDAwKClZWxmwMjDU011u7O5x/fIlJts3wTcIVyNj6oRHwwLrAr5tM1xTYAqDEJrhaJWJ9Xz8k5/mueefxzvHV65c5oG7jjPUEuU9rrXMZjOQAtdaGudomob9yR7bWzeZTPYpBwPMysqR43efe+tke3r3YRG6484fgCiEiLe6FoQs0vbBZ61WgrSkj0gtekp9fqy7SnCwKCznBr1G0fl62HFfq4AdLESx78ASc08So0Ko9Ho64fmoLDB3nTkZbPt/avYn7x6trT545K4zbxmsrh0fDYfIGClNkZ9bkMLjQtYkxUDlGvYmE/b295hUs6ra2316PrO//Lc++PkvfKMs7xuiCCmlpiqqF10I7xZSliEnrAaRlcpR9Fny/XBfyKSOz6rWqDRbuzeZTOtE141w7txpVAj4piXaFhkD2mi0EkTr8QJCkDiXdD1N3VLXnibApAncmOxzZWeXnemcoBTCpPwTZx1aKIaDYdpMvcf5CNGjVSI4eOdo2wbnk97GaJWhhnRzG6VQRZFSW32kbWpaPEpFLt+4ydrKCoSIEZJhYdBCZOq2QJL94ZTECoER6ZQVg6epKwoNPuakSBTaGIrhkGJUIkWCQ9q6IQTBxmiFM5tHePnadRot2ZrscHV3m3tPHyV4QQiCGBTeee6/7wHOnbuP1bV1XBCsbmywtnmE7e0tIg6kYtA4WutwEbRU6CLpOzpJb4InBVpqhIwYI9lYW2FlVKKFZGAUa4UiVjOuvzJlvr+Pq+YMdGINeiJKkq2OHESPMholDREDRYlSBZQDvvT0Jzl//gLettiqYmNU8uC5MxwZDWiqCc5ZZvM5tm0JwWO9pW5bZtMp09kUJRJDsNRGyNIcr/are4FPHVadWzf3XubDch0JS0VIBFLUgQwooRBqsdkHki5uEVaXf/0anctyAVoUv0xmeI3uJ8H6i+8jXqMALQgMXSxFYtMpZZLDARGtPVXbEkUcnLr3nm9tW/utxhiUUhSqkwaI5IwtBD5a8JEQkumud0kWMZvP2J3uh3oy/VIzbX7NOj7xjbS+b4wipPVUefXZNripQm6Q7XlCZqSIPmU19o7QSsqFWFUEopRcvnGTxgek0YTW8S1vexuj4YBoW0y+oQSe4FX6nkLhQqRu2jyjCdgA07rh+t6cq3v7TFqLz6aFIaYM+/FolbXRmEIXTHb3aG1LOS6RsmA2m6VBqhCECCG4pHnIsF0qnsnV22jN4MiRXIQapILdnW2U9nzl5Uvsra+w8qaHKIJEyoiIAh9snp9kex+pCC6glU4Pu/cUWqTCZTSDwYCiLBkOB5SDYXquQuqanIusNJEzR4/x0D338IVLl4lKcPHaqzx671lOjsa42ZxIZDqb8653v4f7778fU5ToqDhy/DibRza5cCHFZmhZMB6PUW2T7Hq6IEIZ+hOlIqWpEiNaRlZHI46ujzm2uoKRgqE2rBWKevsGwaWIbmnbbGiZ/OYEnrZpAIHRBqkKHIagSlQ5JEbFK5ev8fsf/TjDUUkJ2GbOg/fdy5HxkHY+o1CJzNI0DdNqTqEVrW2Yz6fMZjOcc4wHA4xWaAkxio2B0ef+i297vPzZjz/XHJaeA+UhnQ9SitWiOLBgtHa2W6nCZLftmNzyO5c4QrzjyCby2iF1t8JtQshbfn87PXu5oN0JkjtQkIRYev3ZjUMmREMpxaAska2gVJo4GNDUbSJKxECwnmIwSK9JAjbH0IfkGF/NkyNC1dS0VXW+3Zv8dl2Hf/1TH/zs7LAI/XufC71SbRZHX4S4DdyVPOLoi5Baiu6VuRiJnB6azsaSumrY2Z8zrZqkRI5p4I31BNegVZqfROdBWYTQhBBpfEttHbax+CCZVg0396dc35mwXzVYBKgC5zxKGe6/714effgRZpN9XvryCwgR2DyyyRNveQtCCN73/vfR+pZqPidmx27hBd7VSbOidDLYFCJpeKRgc22DBx56kFOnTvGbv/FrbF2/Tl3XiBg5/8olHrz7HKuFQmeXBRkiSiUxJlowECWqMEQfcNYRnUgFriwYDAtG4xGj8QqD0TANdn2CA6XQyKA4eWSNOad4+eZNtidTLl64zLObLzJ49DHWx6vpfZy2PPTwmzhx4jhOKqyLnD19kvsfeIDzF15kb28PITW6UAzbAVVdpddCwtGTFVNn7Q+FKRiPBpw7e4IzR49ybGODcakZmQGllqjsxRd8QPpkyUSU2YVCUJSj1JVGgSxHBFXiUFzfn3H1xk3e//4PsL+7w2SrZXOl5L4Tx7nn1DEKJZChoG0riJHW1uzs77E2HifR4WSfuq4pcsLmaDCkLIdErUaitfe5nXoEHBahAx2KTH72McZlCD0lpS6KT4gBvE/onQctBQSPF6EvHkuh20var68Np8Uo8kEnfZ8ollL1WCZ3H7w6CoJcKm6vOW/KB99kXJr87rSUCGNw3iWrsVIDOUhRdmakC3c87yy2tTRVw97eHrPZnMn+/tXJ1Rv/0jb8o5/6yLOvfKOtr36j3MhSqpsiuKsxxscQt//cnVX7wnxw4SWVnKk1UQhcDDivIAROnDiBgAUdUniUSJ5lMZBICK6msRbrkgh1r6q5ubfP/rymjQIvNE1jUcrwx//4u3nnt7yDEDzv/Tf/hv39fZ58+5P8qR/6IR574i0APPb4E/zcP/h5nL+JCx7nXHfIgwDetxRFgRaCGAWT6ZzNzaMYY3j4TW/iPz3xf+BXf/mXefXCeS5fvwkRTh49hoolAwUyBHwnrFAS7z1BQF03OGuxTYNwAaMURWGSG4MEYzSFKZJwsI+/LhiNCjbXR9Qy8K1veZj505+nsi2f+fwXqPZrvu8938lodcR9m8c4e+5uBqbASYmJHjMoePSRR/jCc5/Jtv0JLnTOU1WKum5SzIKziW4tYVQOOXbsKHedOcXJ48c4cWSDUkm0ACNAR4g2eWgZAR6BMWXKKYoBLUpCCgxCKIU2JWZ1k9nuhKc/+ywfffoZtFK88soF2mnNmY0Bj917jtNHj1AYyXw+QxtFY5P6xHtPVc0ZDEqqumY+T3O98WjEeLzCoDAUhYaiHFijTxglhsDOYek5wEyIQgjfb+x98aGH44KzeGXTPaJUcq32SSxKb0y6cLxIsoYOBTlYHG7rbnpm5VKxugNB4Q/yA93x6/t04kROgOQUbnSKemjblmE5oLWJDSiCo64rlDTJdV9AXVdMJ3PmVc10OmE2m+0023vvs3X4xz/10S988Rtxed8wRUhJta+8vAjUQbASicQ8rAzkgDYBIkRKbSiMScVHBLRRCKEy41Ojle7ILBgpc3wwKZGRdEKzLlA3NbVtaENg3jo8hu3JlP1pjQ0RqTVNG9ncOMJP/MR/xJseeZDxaMhHfv9DXL9xnc3jx/izP/HjPPLwmxiMUizNu7/zu3n1ylV+5Z//Crv7u/mMlYpoCBAQhNYThWM0SCmjddNw7do1trZu8sRbnuSus3fzmU8+zcUXv8IzH/sw519+mYfuuQs9KBEhooRAlxrrHdoU1LNUgLyP1POKtz9yHzKk7J6iNCi1gD4SFCiIKjHTlBGMBprVRnLfiWPsP3IPn/jciyA1L1+9xq//7vv5wR/8k9x18hQ7+zOm1UVMUbAyGrOxsUF57i6+/7u+k89//jlu3LjGjes3GJmC9VGJKQoKJRgMBmysrbG5uZm6oKKgVKlTMzEmUqy3lMl2PHWy0pBY7QK0QQrwIRBl+hmKQYHQBXvTmmeff4H3fejDvHjxZRrraGZzmqrlPW99hAfPHOXY2phCQF1VSBlofWJnySjx3jGZzhiMhuxPJjRtw6AsWVlZYTAoGQ8H6YRdFOXw+PHNatKuHlad22Y1USBsjDGGLEiNMZne9B2RSl28QJLkc51rtUSGJI9A+INQmhTZrkfcESrrmGvdrzIjDOE1Zz28ZmEKGeqX3Rwo3v53QkzPLzIdBoVIHpYiR1UMCkMgpGgXrVLas7VJhB2SF11dWebzit29XfZnU9fuTZ6dXN/9+aiLp79R1/eN0wkpNVdRvehirAVihZwbL8WCOdPNP6WUqQ3uYlZJgWltGwhBJGt475E5TVNrgxS+MwTCOod1nsY6WmexQaAHQ27e2GUyr6i8xaGJHlZXVvmJH/sJvu+7vxulBOfPv8T58+fZ3dtnbXMNG33KKuocDUi+cnXurpQSvfLb54EtMeYQOChUQV1X7O7ucPPmTZyz3P/ggxw5eoTLj1zEqMj5Zz9L1VhGWjEsDNEnGvlodQWlC4YrJaOVFYwSlFpx7Mgmxqjs8puji9MkOLtzp4wdZRSIgNKwNiqJCu49cZyLa6/y8rUJjfXM3Q1+83d/hx/8/u/n5KkTjMuSwmiuhcDG+jrOt0jnue/sWc4eP0rzQI23PlFSM9VbCsGgLDFKE6PPFPsMk4QE0QzKEtfWlIMC7wLW+lR0cwS4KcoEhRDZ2tnmpRe+zBe/9GV29qZs70959coV9qYzgguoCO9+x5t484PnODI0qGDxbUOILSJ4pDKYmDRizjnmTc1sPqeqG4RQDAYDBoMSY4r8+gFjtFFyUGh1WITu0CAE59vgXFgw4mLatKOHqPs8rd4Rv2OgiQ7liETu3H0sD4ruzJK73U3736Gg8trkuSSmpU99ThlmnVZRZJNTERduERFJ8I4gkqxgNm+Yz2uqqsbP55e0ix9EF5/8nz76bDgsQv+hb2Qp5xL5ZUKYgjrWg3CZIpwWPy2wyqaUopt8Ro8xA5SSmEITlaK1FpSkHBbMt/ZRBpRRydzUJzse2ybLnSAFrQvsT2fUrUWbEtt6VlfX+M7v/B7e9e3fxsb6BtVsiq3bpLUhsrW9zQc//GFMOeah+x9BKc0Xnv8in/v8F3DOp2JpigQZOtdrEDypo3Mha2WUxDnLdDalqipiFJw9ezcbK6v4ek6o5oTgsCGgnCUlARuENtgQ+fKLF7Bty7Ejm7hqTlkYTA7ikjqPfTuIIh58dI0xFGVBiMkF/Nh4xINnT3Fze07lPPPZjFdeeYUPfuiDbKytcO7kMQam4NjRo+zcvIkUkYEwqPEYsbKCkhJbVyit8S7ph6IPGKPxrkXJMmmHlKR1jqAMsqDfmNoY0MMBgxWDQ2CtI0TB9t4+06ri6vVrvPDCC1y7cZ2vvPQy8/kcEFgbWB8WnL3rGJsrQ77l0fs5ujZCY/F1Swwpv0gp2XuZgcI6R9NaZnXFvGnQOX69KAoKY1BSYXSy2i+1LAotD4vQrQdIIZyWoooxBu8TxOl9IuIEtWDIEQJBhD5ITvqk6SLHdt9KQEjRDiqnqS5sexZFSNySP/ba0FvMXydieM3i08+IXkvUmhENcQuzrnMDycEMyY6oL5rpQBxwzKc1jXXs7e1TV/OrblZ9cLo3/9Wf/vgL+9/I6/uGKUJX9l62R8tjl7xzu7JIimnRO9wmz6bOJ07r5LqbrNbTrWDbBiUDEo/1nmI4wMdI3bZIrfAq28HnNFNrk8peSomSmmADs2pO3TagBxSDASdPnuAHfuD7ufvuu8F7bNNSz6dUsxlVXVG3FR/7xCc4duwUxzZPECM888wnefbZz2OtoxwOqeoqdR5LgVzd/CS1/+nWbZuGuqqzO0ES0a5tbPD2d7yD3auXeP7TTxOioLWe0WiEGZTULjl8f+rTn6K2sLa6xs3pFCUDzreEUCDlKFniS9HHpvfBf4A2KV5YK8vQaFZLwz2nTnFja5/nXr6GQLG+vsbzzz/HQ/ecoZ3cw5G1dYiRI+sbCCkYj0a0rUIqgZGKWgqUEDidfJCEgcJonEtJq12YHwKCkihtaOsaM17NtVLS+EQ4aV1ga2+PL3/lK1y9fp0XXvgSL754Hm0ETe2p68DICAYicmZzlW9766Pce9cJZHSo2IK3+OgQIqILhbYKX3uEDygkFnDOU9sW6x3GDFFaHxhqK60ISedktJLjw7Jz+3xfwCwGbzvLIx8CKqSCsyhCCWr1QSYuHfmZUB3UcZDx1m/04tb4h4Nfsxx2d2sRey0o7vbu5+uYO/HaxYmlZ6qzFuqhyJD2m6pNeUO1dbu+aj40nzT/0KM//42+uPoNdjPfjM6/GkN4DCmKvLQpzTAuiAhKSJSQ2cInuWiPhmNKrZAyMhwMme5PsN5CUSCMIuBxWa1v2+QJJ4TCaIFSBV6AEgYhEvHp+77ve3nXe76L++6/j4CntQ0Bh/eB4APDogApuXbpKr/wD/9//MOf+4UkgPVpqC4luLZlWKRBeswzmfRQpYdGC9AKSqNxOYtIZu2TtQGpYHVtjR/54R+mjJZLr1xAxoA0BbIYYozmxv6EaVWzN50z1DVHj25ydPMIRZFp0SLRTGWOTE/qdJkx+IjQCmMKvHOUpaNsJaeOrPG2xx5mNF7lCy9d4PorV9AKPvXJp/n9D3wIb9Mp97/6L/+PDAYl9913Dxtr6zSzmmFZYl1kZTQixIrhoKSua+ZtYuQRA6aUiCBhlBwxJtMZEcmsagg+8NKFC1y/eYMrV67x0Y99gnlt08mZQDVP76+v0t61buCh+07z9jc/wb1nz1IqgQxNPnBIbPI56u+VbtMySuN9RKGwwdO2aWieGIzJtLXbjLRQ+HTONUqIwWHNua09cG3d7hS6bGMuOssCU5+9FcHjhQSZoWuRipOUPpkHd91ISIfDlGOZSDghExa67ufWsLoouo5K3N4BdZEod3DeXi46iz9fGPfIg+onJGEZnMust3x3dT93yEy47MLvnaOqW6bTmu3dvabanz1V78z+NxfVx/7Ox591h0XoG4mcoNWeqMOzPrhvV9IcjSLRcSU5oySF6yDRkC1ryKwpJeH06ePsti3Xd6e0TWA0GqK1IDidb7jE77fBE6NAG40qFEEYdvb2GI9GzK2nWFnh7Lm7eeItT2BKnTN9LN61tG2dikUEow3WBebTKVoXPRvIGI3wyUsuxJQuqVXnRh3Bp83OFAXGGAZliSgLhuUgFdcQsdZihCJEjylK3vmu7+D3f2/OfD5ndXWVYjhiuLLC+Wuf5eGH38SL588z3Znxlsce5ejGEWK9m2Zoyw9qyLBB/7BKRBQU5Tg7TzhKIwmF4K7jmxzZ2ODtb3mcmWv5rd/5fV5+eQsFbG4MOXb0JL/zu+/n8rUrXNvewxA5e+YE3/1d7wHgrjNnWFlZoa1rirJESkld11x69VXqtmVQDlld3+QrL7/Mv/j13yQ/t2gNKysFUkom+xPqJtA6KBa5Ytx/+ihPPPYg9959F6dPHGOlLFPMcjVjpA2+DbiQcpEKVeBV6pBDkEhhEaJNOWX5fbDO0rSKKCQq2wul1F6RZ3qdHCAWSnLYCd3aScRoq6ra1wPVxriIcPAqIH3Ae4mXOlOzA1FCkOnXeKsbQoyQ009v7Spu7V66DymSWeod4bilbkhkFOBW2vet3U+SBx1Mv3tNi59IsovK3V76+ZN9l3M2z6ot82rO/v4MW80v7t/Y+idI/YG/+4lnvynSfN9QRchouaek+pBz/se0KY4uqNiBmJk2sdtYU/9LVElDYtuGUidqtnUeYyTnX77IH3viMSpbEb1LztYx4LLyeVCWmIHGC83aSmRWe1Qx5F3f8308+bYnEVLQ5llOjBEXI8PhgLX1VcqyJITIqCyROedHKZVseILHqFRwtFIUWvZGpjFGUJGyKFgdD1ldGWEiKK0pC531KUOUBKM0WEtVVdy4cYPxyhrHjh2j9QFdDrh4+Sr/6nffD0oym80wxrCyukpVzRjIiDEGbUzyxwsxwVIhETRsTD5pzsUUWSwNxaCktAXWWVRTMxKa6ByDQcn3fsdb8Erx6Wef5cKFLXb2LlIMblDZGoxiZWOdSYg8+9J5AF589VXapkFJhW1bnPdEoG0s1lnaNpEC9vcntLbF+7RJWB/ZmzWYbE7rA6wPDPfefZZv/5a3c2JjHUVkfWXIuJAUImKbGSo6ylIihaN2NdElI1RQSE8O00tdDkribYvI2UPeJ9hEaYUUidUkMtMqNeEBqQxKCGO0Wvkf/8x75H//6x8Kh+UnXT//6S/Fv/zImV0lxHx5JiT8Ihco9POgkCBa7/BSQNBIF1Gqqz+yLz5dJxTj4jN3pk6LWzoZQKpFUXvNYhO/OjlBZMfKOxStuITMpNyhnPuV/fG8d9jWYl1NU1XMJnOq6WTiZ81ToD/ydz/x3DdNUOIbqghd2rvijgw3v2JDeyHi75dI3dl6SFJWvcgtbyDi80lEEJF4NtbHjIaGjbUBG5snePqZT3LPiZOc2FjFVgHv2nx6SVCXKQzlYEhAc2TNMBiMkaMxf+zJN3P36TM0bYvSJiUtKsHKygrrmxusra0yGo1SxLd1yIGkaR0hBFZXV/ND55IeAoGPDkWy8AiZnTYcFKytjFgdjSm1RmQG2cpwwNqwYG93m62tir2t68y2ruPrGceOHaNpGszI8Lnnv8Sv/uZvceLECS5cuMDJI0e5/6672RiXEAMroxW0SpZHWggEIWX2OIvA44LDBoeMmugCzlukVChlWBmP0MIwn9VoqZi7hhNrY1Y2j3DiyBH23l6xv9ewtbPHJz77OZq2ZXv7JiujEZ/97A4QaOuG4XBICCkLSEqJtRalVOp6YipIUiRDx0ImUOPu0ye4//4HUFJwdHOTtdU1hoVhdVhyfHODImRn8eCJbc28nqVjSvRY12Jti1QK37bYNlF+nUvWSZZwAHLzLhKlAAciSoxUaU7lbSKfSEFAY31LoQ1SllopNRbCa6A9LD/LKEaxLbXeb52n8AmWlgFCUPngF5LGLWQjX5HEn5DCH9O6eEJQiFxA0iEkLIFfyYdQynig4Cw7G4glceqdio/4OmZEXxV5vMXXLpGmfDZpzR8+JOKTbWmyP+S8qnxoms9OdvZ/MYjiwjfT2r7RZkIMiuJ6O6+fjq17R9T6qJQynTLEAtPvNdUyt84+IrCMjWRtZJg0iihga2/Czb0Zp46fRLUt0jka22A0KC0phgOEKlFSMYgCaTxHjm+wPjDE2R4+SlaPHKexLs9OSopiwOaRo5SDUTK4LIsUymZSxF6IEakMWpucHBwxQkOMGJmYM8F7VgcDNldWGGqDVprBcMzmeI0Vo2n2t7GTLex8xnzrKrQNRqbhrTYFV25s8+JLF7ExdThhPuXk3ac4e3SNoY6USuJ9QIoyWxt5XDtH5VlQ9AkukSHgnE1WJNERXKBQBY3zgE2svTZZHiljMK7l7OoKJ1dGTEYVe+slk93jVDFkj7lUcISUqPW1ZGEkJXowSp2kSZv/YDBAi+TFVWiFbx1CClZXR5w4doxzd51kNCw5srHB6niUmH4CCCnV0jdNJjhYrEsdlQ8uCx2hbmq883jn+xmQj4HgQUqN9PkkqyC0AekF2NjPJQqtETEF8ElA6FScXLBlFHEFxGERunVzVno7eLakklGIKCSOICJOBBwFOkDEg0/PZhAQRLazzdlCREnSvMpFcnIXxy1l3yUtdyW9QwLJtb0XrC5/3VI341lY+/RzK1KEiBCiz0ISKCIBj+8gx1QwhcpjgM5+yCeZQTY0jSF14B3937b5o24vV/uzX3VCfeR/furz7rAIfQNfl/eu7R4drL/fhvhjII6GjpQQuxswhcdFIVA5obEbFmoVuevkMSob+NLLr6JUyYVXLnPXmTNslEOaZs5otIq1NeVgkJwLijRnLkYlUQrK0rB99VW2rt9ADkcMtaEcryQ3bAXHNte5955zXLt6mZcvJrp2MSwYZIV39GERS5xxZSUybTPPrgZmyOb6OsePbGTorWA0GnP/3WcJ9YQrV3bZ3b1JdC3jwRAfDUiJ1gUXXzrPJ575FB9/5lN853d/D7/xz3+J1cJwdG3M8Y0xRkCwNZhhso1HEBpLqxySBI1E51OGT/B5pBr7DlEE0MIwKCJSSIrCMKsqqnqGdQ7tA7rQnNgYcfrEBm9604OY4QjvArN5mllJnRwptnd2sNb2p9EQAoPBgLXxiMFggDGGtdXVXlisjEILgRKRtq5S2KCtidHROJvcF6zF2zTwdc7ifMB5l4fCIZNDEhzUrUN3OvZhcTJWpHiLmC1jYhT9OFrkTYXMhuoynAhCC6EG4MRh2bm1FTIzEbjivK2j18PYJZYi+04o+kDE4rNf3ILRFhA+SRWWPeAkqWAJKV5zJvRacNqdIbb4B/o7t/MvcicUYi4+HlxCPdLhLuDzh3NZg+g9rfPB4D/nbPyd//mp57/p3Db0G/F+Hg9GL+w08+e8D/cKIYZSigTJxUhgscmD6PNJCBE1KDl59Bg7+w0vyy0efvxNPPXMJ7n3nnOs3HuWYnWDZm8LJQtWx6sMyyLrZwJlkRXXwXLz6mXaAGU5JtQNg7UVVlbXGI7GnFxfobnrLJe+vMHe5ZfBaHRRUHufNEc22dZ3V6KAyxzHAMOiYG1tlWNHj7KxsU5ZGDY21okh4Ks9Ln1lhpaC9cEQGOKERBUDnIcvXHyJf/m7v8uF86/yIz/yZ/g7f/9nOTUa8H3f+U6Oro3ANcxtw7goWB2VGK3w1uIFRBcXw9MQEblzSYwjn4kBsScvKCUY6ZK2bQm+yDHNHttWVI1HCp2IFXqCKwcYU7KmNRsrI3RhMLrkrrXVPlsmqbw8SqrUnUmBj1C3yZDVti02O38H71IBihEFONti2wbvbOrcctFZHmov7glyASGn7oLMlGuVOyWBwEoJPvR+ZSEEtBa3QC2xP1KnoDahEaKIURwWoVsvqaoYuUmg9iEOpcv9Yj4QxOhwvXuIzM7U2RBUyJQvFBYpqVIkpmu6fxRyiWfQF4wYiR2LLs+OUzQ4rz3reQ2OtYh3/lxvnpz/PbF0z/Uz6hARPqcr+3T/tm1DVTfMm4b5/uSy35s+7eHiN+PSviGL0OqwvDmvq/dNrX+nLOTdXTudNoWIkiKZd3aDwRiQKokiSyO56+RJGqf5/Oc+z+OPPsGv/dZv80N/4rv5liceT5Y/IjIeFti2RqjIYDBIg2mlkUrjIgwyJLN94zJiR2N0iQs+neCHJY89dD9HV4ZMJ1PaaJFGpvA4n1JVl09rm+ubrKysIEUiIIyGBUVRImVEkzBFIUOKbSgHqeuTiigUbVNz+cYNXrpwgfd/4AOYsuDUqVP8g5/7OU6NRvzg976LU8dXEK7GtzWllIwK3ac3CgHBtgu8OqR0VZkfeBdtMpZk4fnVm/SJZNi4Mh5SFAXTak7TtEl0iKf1liBqfDPHSo3JwlwXPFIofKbTC60YKIPSyaEhUVdTgmnIp13vkpYn+uTHpYXEujYr7X0/t0odTnrYE5Mt2+XnmA2RIZ4OqumKUDKSdEmc2jQIkXUhMtOCY0AIfaAAxeUNKMkUVUSUEeRh1bm1SxA2xngtEufBh80QBNILohcEF/DK40mQFzImckKmQwsRETEgolysmxTp93mWuoDeDtKz42vMbF6Lio24fbazHJx3a4HJU6Sl+U+KGw/dr/0cKBWf6Cy2banrhqppmU6n+5OtrY+FJv7L/88nvzI9LELfJNdzVy7UD26efqquphdj9GeUVErluG+CT5HVsts4OpVyitgO1rKiDQ+cPsWrr1zm+S8+B1pzeWuH85ev8sjddzEwAiNTHpEuEi03BFC6xBiDCxGkQkhJiBFTlhAlpZYIAto6joxGrN5zT8aVHcg+ECWpwLMSPLGvkv271im0TetkZSOyo7TSAqUUtnGE4PBBU1cNFy5f5gsvfJnf/K1/xV/83/0nXL5yjf3dbTZXxnzPu9/Fow/cTyEcfraF9xUFivGwZFQaVAwE55Ay0mZoKiwrvWMXwXyQ6RN9ghlCdgn2EbTWDExBWazhXKBpG+qmpWkanHcYIyFaqlmFDwvle902SCRCSeZaoZW+bVAcYprD9B1N9FhncUrhvU3ZUCKdiGWUIEGTZjQp2DAXIZFjokV6L3uW1ZKtio1pHnebKl+krrDLs+mLzq2UXNA+xjLEwyJ0hyLkqrq5JKOcuVGJjiIz4ZbWlpAE4vFg6F33DEtxEC4TiNv0QGRNUMy0bHFLoelnSbeWp6+jd11eexH9AW3iIiHWJSf3TECI3qdEXuuIwePalraqaVtL1TSuns2+GCz/KEj92W/WtdVv1Jt6c1huTar9TzsR37w6LNeJnmZe422TZ0ARHxxBBZQA7wOFUXgPY6OJMXLfXWeoXnmZaAZcvnSF+WTKyaPHWD12DKlhMBqhdWTe1JTlOG08OXZYStUPQ7VSOGeRyuC9x7UOJSVDo1MB8xZwCBn7EPJkE5LYP7KUSCWyyWog+OzfplViibUtEYfSBdOq5uq1a3zu2ee4sb3HyVOnMEbzmWc+SbW3y5HxkDc/8gBPPHCOUQHtbI6RaWZmhMIogVEqkxMszvoEYSIQIvmgCZJTg5Qqx5unzT+EgJeS4AQRR/AeKWS2OPIURZESY5VkYAxGa5rMeLPW5o3B09Q2x3CALnQ6wSqV/bYWEIaUaeNJkGDMgt5k8W+0IupkvNoVFJVp70oplFTZuinpRKSQaC072GxhwxI8zrocIbBgUCmlwNulrwu3ZdZ0BWzpxK1CpIiLAeXhla9/8MnP+f/sifuvGy1mLgRsiOggUEGnMDuybqiDTvvuRtwxklsKmaG4W/OC/mBpql+74Nz++eU014zCZfKBT15xS38eQpI4hOAJ1uJbi3Up2LGdz16x0+pXvdAf/XtPfbE9LELfRNd/+m1/TFy+uhW3fHstKlMf3xitixjZcTWzapIsfEQarKPSXMgok6zhvUPQMioHPHjPaa7v3WS/adm6cZWmnvPcCy8wKEtOHtlEm4JgBKUuMLrsb75CJJFif1LO3ZBWihCTIWhn0igIKco6M+A6n7YoVcq/6U5vIc0XpNIImZJWtTLUtsF5ydWtbS5ceIX9uma0tsZHP/UZdnd2eMfb3srIGF78wmd55Owpzp05yX3nznDPiVVuXL9KbKc09YxxWTAelwzLAhEiTdMkw9bcIUipUDp5oaU+TWKUIkpwJNPPEDw6Juacsw7vE3SVyAUgPYyKFYqixHmHdYEiRpxPHCItdZrhhDlSQFmWiaWnVHYVpof6usG1yqdZrU1vZdQVBKkkKhdJKTvoRvSHg+QhKHoXZSVTi9INkEMIWBtAJeixtXl8QbJRWr5CNqC9bWM7IHyUMgphQhpVHV63XC6KLRXZakPEhKSdiz6APjhHORjXfQfCgUwf6aAklgqW7GNcX9MlW3azQflVC9BiBnRwtij67KNbEIK+E7IJcvdJG+RDuv+dTUXIWof1jno+351u7/xu24pf+Zmnv3Tzm3ld3zBF6P/1l/9cGZw/UlfNeHtnsnYzzs8qax/WsRVHh+nULeoBotaUOuXPyC7iAbDWIbRAK5Ow59iyvlLy7U8+zsc+87l0so6RD3zwQzjnOHfmLE888SgbgxV0MSB4m3zUhEiuyQS0EGitCN5l+mdAhJjTPSUu+F5hTxa1+ghCJm1R6j5S4ekBhmzJM61rtraucWNrmyvXb7K9v88HPvwRzr/8Mj/0Z36YlfVV9vd2+MB738taOeT7v/PbefyB+zEqIkLD9tVXcXVF8A0r4wGFNhRGI1XqrrpYcaEEUkuU0snZWpnFHEWqNBPJ+LbMNPjoU3Sxdy1aFxhTUFWJ+da2jvWNDQbDISaC80nI2dYtjbcJthwMEaQNI23umZbgfSJF5I1GIVLUundobfquRy3BaiEkeyEp5cJOR6SoAJm7oN5DTMReB+K9p23bA6r6rqPqI6eXNCWdg8JCCLBAcRYncSFBmBgPO6E771ZmW0le9s7XzoiB8jLHGETI2p4OjhNfxQGh74TEIol42R+uJxl8FbbbsrC1Mw6+8+zo9r93e5cU+9lz8D454AfSYc15nLXpV2epnKVqPW1TfwXLr4F66Zt+Wd8I9+7P/Td/6e5zd538z8tSP+4jm23rVk6dXbf1Bz58qo1q7ejIMB6vMFKRjVIyGgzQkDn5iQWllSFEUAKkjNTtlFJHTm6MeM+3PsnHnvkMFy7fYLA+5sbeLr/7wQ/y4z/257j/7F2MhoZjG+usr44oBgOct5SmSBuQEslyJ2uSQi5CkYhwILRO1N+yTLCXjxiTXalbj1IaGwJV01BVNXt7e8QIN25e59f+xa/xmS+8wNkzZ3jiLW/hPd/13ez91m/yW7/+26ytjji5ucJP/Jk/xVsfeZihBDefMJ3s0VRTXN3gbIOSgkE5YDweM9CGtmlpXbIJMkWB1BplDMokiyClEoSoM9yIygEZveVI2sC9c4RQJgJAbdAmRZfv7u4TpWbkI6srKwzKIRHJwAzwIRcGrRAoXAzppJhDvhBLRq4iG0/K2A+Gu9Ouyt2jJHnLyaxcFxkbSUy+0JeLzp9MLsUFxBj7jilpzfwC6lkucq3trZZ8CIn2L2V2Soj9e5I62Sh8jCrEeMiOu8MlpNo3Rl2qna180AMXAtpDcJEgA0ILQvDIpUZSLMFyiw5X9XO9ZUhuOR/11ojvRUsbc38TbilyWQDbER6X5pDLHZD3bsloOPZecLGLpwhZ2iBSRIO3FutTB1S3jnlr2dvbvx7mzfs9+pM/8/Tz4bAIfYNfP/tf/sf3bawP/7u9avbuWIWTQsqVcjgqH37sYXnk5DG2d/aYVw2NC5jokbbCGIUUIVMo0xAy5Na+604KLVHCYXCsF5J3PPEYZ87u88yzL/CB3/sI3/297+aLL77ARz70EaSI/OgP/ykQnuFgwOrqCpvrqwzLktXVVWzTYLRJiaw+gMsnbATBOVyAgMNlQeRkukUIgaZpEVKzP9nj5vYOL198mU984ila2/Id73oXDz72OK0QXHz1Ek898wlCaxEIfuh7/jhvfuwRVgaGE5vrNLMJ87ammk6oZvt4mzbOski5N8PhEGKkqmuCTxupKgrMYIAyBTrb92hj0CpDcl0RWiIKdPHL3lu8lPigsvVNgvTatgWlmM/nWJtiGtbWFEZLdFHkwqJSN0aO4g5pXtelZfYn2ggoiDlqQsQF+iVC0ljJ7hNZw9THAYRI6HJdlpiIXdzH8kl5AfuIW0kGmanVsePSvdPNspZfawcP5bZbHHZCd76CkM1sVr+sxmoSYLMr3iE7JfgIUorbMoFunfu8NoyW/FNEBpS7LluwYMkppV6zM+q+x3J3090/xHiHzqqLofBJ++Md3tkkyg6uF0l776maiqq1TOZN5ebVx2b7za/8f5/58vXXRYP7er5p//Zf/DNHBoX8b6oQ/6Sdze4dlxqlJG66x2i8wj0nj3NkZcxkWjGtai55i60HqTV2jqBlYsEE0jwgs9kIPs2MnCNQM9IDjo2HrK6sEAg8/fmX+NxnPoXzkVE54k0PPYKXmo989ONcvnyZ4ANPvvXNPP7444xGI0bDUVJBZyGqNrr3lxJC0tiWpqkQSvH881/kE08/lZgzCDaPHOHRxx6lNANu7O4RleLSqzf4wEc+zGg4YG93nzOnjvHAPecYas09Z05z16njDI0C1+Imu8yn+9impq5m+OAxSqO1YFgMGY4GaC2om4pgkwu3KQcJLjMlsjCYokDr1M0opVOhyJBcAHynnwkRhEN2jNUgOr0mKkSUSXOx6XTK/nRCWZYMigJZxmQR1EEoUiIFyCiRZe4a00glz2KS62OQgiB0z3KKWYneaTFkzhhKJ1KJiMl/TIiIEj7j9qKHXjrK79c9nF6CZoJfyr3pilhH4b4FOYrxsODc6fqFT33e/oVH779QmLBrfHlOA9FHhI55I3cIqW+JY5AHOtbeFUEc9Hjr/w49/TKxIZEH1jIsG6HGJUw1Ox90xMYYF04IMcZFDENnStoLntNrd96mjt6lw26wFu8s1lqqumHWtMxby3w2v1hP2l+Isvj06wZlfT3ftPVs71vjqbXvsnV976hUBNegVIFEIL1Fac3KYEChC8qiZHtnFyUVzrt840AIAqHSZpFglIiLAQXIDC1pFVgZFlBbHr7rLGtrK2ztVzzzqc8xmc05/xXB9t42r7xymfl8xtr6GrvTilevXmdz8whm2rC7u8Pe3n5vFEqeF62urDIYFjhb0zrL7v4ebduyu7tD3Xhubt1kf38XrTT1vGI+n1JIWF8d8cB997C+tsrJo0e468QJhHNsro5R3mPnE7x37O3t0toa6z0+pNlUYQaUZclQD1BG0LYVzlqi8xSjgrIsMUWJ0hplNErrBMtp03cpfRol3QE/5twWcQDyCD7NiyAglUTr9P7P5zMaWxFYJeD7E6UPyd1cZEEqJA82Seo6upMritTN5N+nVyCWTqZkx29ydGfyC+wdHohLxpa3antuxfXvXJg6Gm8/F8u6ICHvzNpKUGUQMYRDOO61uiHkxejsq875N/sYhVcKML1+TIREIPlqpIF+/cPinuziHW6D3xZ9bV6jcPvch2U9Ubjl37kDaSKE3nEjLAm8Q0wyh+hyKKa11E1D1dTU1lE17c3Y+t8Jsnj6733i2fawCH2DX3/1h7/rRBuaPzmtqnsHClxI9vkNDmMMPoAJkcGgRHnwUbC2ssJNvZWySTJmHGJAY3L+e77hPAid9DhKqgTbOMdQS0plOHX8AebW4af7NNazP2uYbt9kZ3ePkZFEb7l66TLBOV4tLtO2LXt7e8zmc5q6RmudNiolGQ6GjAYlg4FBCJhMJhAcWgiMgBVjiPUcYTRHV4ac2hgzfmDAY489yrlz51gdlYzKglII2vkM38yYTvZp5hVCBHxbE4NDiaRjSjEDhtFwRKE0zlvqusY5i5EKY0z60BqZA+u6OZBQWQRIRITlzTl9LnI7VJG6Tp+92TzISAgOZxucdYkZFAO+p10nY1kZu+8f8vk12yRnxl6HZ8kYU4Bh6E6vYgkaSfBNyPHPC4J32hSiSCmY0cd+VhSjJEZ30GgSQUAezJ5Zmit08GDnkCByHHoHVx44jcd0HZab15wL3TSET8fg3hWk3OgslJSSPeMsZOZiF27YzQgji4C6kDBZ8EnMeqAbEksC4w5+Rd123BBLOF5vg5oPObIrQLd0WgeLUkhShdiJUUNigrYuzUydpWkq6ralbd3cz+YfsXX45YC89Hpa09dvJxTsfStH15+cTfeOSC2pg2M43gAtKWyarQQPY6XRekBZRMajMWVR0tQtUiTBovcBL3waegrQQqEC4CVRKWJUOd3RoZVEE1HVjM3hkB/7E99H0Jp549ja2uFDH3kqOb7IyHS2y8UXbuCDSAr7THMOMeKVyHqFSLUr2PIp8kxKzerqCqc3NgirGwwGBY8+8iCnT59mVBZsbqyxMhpR6LQhT6f72CYVnt26wtZNsqixDa61eeNPxIsi5w4ppTHaMBqkgLiqrrG2JYqI0gq99KG0Sm4B3UyDjh6bYAuZNU39g+c9MSTY0fv0oHmXjUJtUoLbpsW7pmcDOevw2icNiFH5BJszVmJyoSCkTT2ktiOxR7phcC6I3Sk069PzCTjgPUsRHiBkzGaVkui62PeF9X+MaSTdkUjCEt32wP+LZL2/yK3JwsmleZBUsjtfd/b8McbolicLh9dtZWhSz9tnB0W84dWoL0J4iVAeHyUyyETqWS7waUTYHwyCCP0s8mCnkhzTl8Wry3CckPJrQq9dP7RMwabrrJe6n64b6pKYrfVYF3DWEnK+mG2rlJq6v/slu29/2Ynysz/z9BfCYRH6Br/+7z/wx0Vw9T1Vo85EawGLD7Azs4xXVxiWJQiJVAZZWcxAETxoaSiMWbLeSGf4kAfPKbMElNAQJM6CMAKlJdF7CIFCCtrJHitGIW1F7SJjU7B5ZpPH/9KfRqCY1y2TqqZuW4RSbN3cIeZBvo8BrZLbQTfcDjEghWJtdZUzp0+jlUEQUUqmHTkGgrUE1zK/uU8tIsE6bNMQY2TWVHnYmYwerbPphKgMK4MhMkbKwrA6HidBZgSpRXItqGfUzRytFbEoMpsob8bBp5MkEH0HWohcFCIhz7WCS5XDd6QE77C2xTtLcJ6mbbFNQ1PVVLMptm2AZJ8jokAEgYwiz3Cys0EQPadAqK4L4QCJQMQAwvfiVZYGxSLrN0JMHU/XDXWQiFjWbuRNJmRzyRDB5fwnHxezph7Mu4WwEGIanEu/2ARlpt53bgqBgA/eRe/qGHGHxebO1y8+90X3Ew+cfZ79/ZfKwtwbhDHO+ySAzum+IgqiCIvRTZ7xRCJa67zGycanZ6eJeACqy1RJ6IuOy93R1yfhyva0S4XI5wNUeg6cc8mj0Ht8SOF01iYRqm1bomto2zqRpqr6Sn1z5zeiWn3/3//0FyavtzV9XRYhb9uR1v5cVVWbKkJVzahbi5NTxvMpg2LA+toam5ub2BAY5LZdypiYcTLZyXRYrydrcrr2WpBjrQNk94Oo0im7bhqUklTVDJylWBkR6hlOKgpCsutxjuNrIyJjfAycPbqZ2VjpMoVJG2LIlOD8OqRQiGCx9TzPrmyaXwWfxKPeE71DCoG3Lc657I1GCn8LKfitC9yTQlNoxWg4YGAMg0GREIquULg200MtIHABWhew1hGFRuKQIaIMyJjo42kY271zorcgIcTc3bR9ForvkiFtg2sb9mczprM5jetiD3QP5oUYEd6nJFyZDCmJKRROiYiXKndeiQDhY6qMStLrlGIPj7AABzMhIfkHdkuaWVd5sTvYsC800SWLp+ggOmJ0ucbFpX8js+nCUreTIT2vJaHTpsRFxHOIwbat3YvxMMbhq/ZCynzFN/MPedu8zSpxwgSNCQpnk4u8xyNkJMj0PocgiC6LutVBMatY6oD6GeBS9yPCLdZKItzS/iz9uRB0vvGih+T6gR9EegJSXD6QZQKCaxts0+SwOsesadmr/azdqz4QxPA3f+bTL155Pa7n67IIBWsNKh4vi3LgnMXrEtsk+uPe7i4zpWltQxSRTSJSCbQxROHQJgkPfQ8rpQ3Ly4jWMm+sHiFDTsmMeJ/uWx8CUSbYLvqAEg4/nSGVJGpDHasMBQjqqUWINFwXqoWc7Arg2oWtSLd5+hho/VJh8mExrM9tvXMJ4op0Ds8CH0CpxBBTOukjtDYURTI5VUoyLEvKQqOUIMRkT+yDx3ZwQQDhA03b0rSOovBE5dDCpCIHSNdltXBgBrI8fO2GrW0HvbkW5yxt2+KsZXdvn1nd4r1A6xKli+zllYp9Ol36ZOSamXVSSGKQyb0hG1CGTtSby/dyFhDIBbEpZPbS0rwqFVCVYDwREj2f0M9youisVVLYGCEHjnWQi+ggORApywGV+rp07wiISiN0nqNldb2NHhtUW7duOwgzPyw1r3390gsXpv/R/cc+7V1z2Xp5wnmJMUXe9mVynZY5jFKkz3aR2KLHVmNfGIgyuaHEkBlxy9PM7rCSNGXittC5pSIkBZ6AJwlmpUgdfBbKJcTCu/xa0n7kQjqQOdsQXQtthWscMxfZb6Kfz90nQy3+oSrGn369rufrcyYUghBCDrQxupsb6MIQbIuIEucc08m0F63pwlCSbGWkSFg90aczuFDcwsVkyYJy6Yak51WlPBDXxwcLIQgmDR+FVOmGFKrnj0mpkp9uRyXuB6iLLsD5zN2KaTPrs+bhYPZ8N5PoqagSqRI1XalELCjLYU8wUEoxKDQdszkN3Q9aj6QMkxYhJKORTZoMvyg4wiVWXd9NLPmlhZCEqd77bD+SilDbpCLU2jYVIedomjZ/X4ExiXlHLqYdDyFREXI3EtN7FkiarrQGYjEQTi8iJ+RGYhALbJ7MjgqJiLB8oo3ZCZwMwd3qet3BdOIAdrP05xmG7BJZffR9fpAAtEiC2WBdFt4KnA003rVS6q3ohT8sNV+rHTLPN5PZM8VwcL/zYc05x7AYJQhXJ5EyMhBkOkAECYjQHxhEv365QIh0QBGRXieUaNcq0bZDPgyFeEdqd3eAiTmlOUa5kLMu3TMxJvKB6wITs0NC6wK+dVjnaYJn3nqauj1vp80vajP8xN976nPhsAh9U92gwglEo5XyoiiS55hSVPWMECJNVVPXdR87gBCsrq0RSGI0rRStc3nXi/2hKSUfxv5g1OXhpUKS5x/d0DH4zM5JG2VrJSbHASyLG0PeSK31yf16iSbai9uEQOW4gOUN3rlF7s2yIC91O8lGRwiBMQatNcakDsiYAcZ0f57m+JBOacIvVN+dFY0U0FpHVVXM5/Ok/s9WQyJb5yjVWdbEDGGlDTh4n+znMw7e2d00TYNtmxTKZRNEN5+nBmA4HDIajRgOBqmLlDIV6SiXiku2wpeZBh6yJdAtYkDPghodvEfGg87eCV2JvZo15g4qRSrL3lCyj1fO84RE6yV/dILJ5KwQ8q82pAIUMulBRjARVIzoSEqz7dzHhSR6vx9CvPi33/vRcFhlvhYkp6408/DbKz788cb5NWMC3jm0STdEcsJWuTsNyZFEZOYjPvfIGWrF9/lDMUOzHdSWDn0BEdNhZzFkut2kNM0uF07ykYR6RBaElRgizjsam2I/vA201tM2gabx1LVl1lrmVXPdTerflEL/m5956nN7r+e1fF0WISF1G2Pc0Uo3hTFjQqAsCgZlkfJeTEFd14kavbvXxyEUwwGIiFayT2yk3/RFpmzmyUOXIaxSQTCFTumZuRB4F3oTUvLp3TmXWFcx9ht493ecC70VTD+w7plVIJzri0v3NcsFyxiz8D+Tsi84Uqb0UqUVRhe5IJmlKONAcL5XixOXXbDT9ysKk7PsW/b3JSGE7Hit++LbkQRCP0/p7OgzC847vAs5sdRlCMISgSZ3QzFGhsMh62trrK2vU5ZJiyRVgll6a/3Q95z4YA+4WiPkgSLEcoxzzEy5roPLhZa+e6UnLaS5ge8LVpc/JyJLUONiY/HZucGHmNY+Q6ghl80kgE2HFY1Ai5T+GXw6sNRRsLW1tT2d168clpivg6DwwqvNX3jo9Keaaf1UsV7cFSMrzrUUyuQUW42ICQ5L8xmx6HASELGA5SSZOZnpBMsBhpms0q95tm4SfXdzAI2jGxl1sHunFYgiUb6dS+a9TZNYp74NtE1L07RUdc3cWqrG7rpZ/V7bhF/+uc8895XX+1q+LouQ1NoKGXaKomiM0YhM4yzLIs0lBgPqumY6mTKv5kwmE4RUjDO8lRx2ycPt7B0mYu9dJrLz8nLi5rL7chK+pc0WFw+kdC4ndPY5J1KiBkV/upK3GCqGvMt3cJrO84TlgtX9viscXecjpaIoVHaM1kvFr3s9C4BRRLLoU+JJIlOtdIop1zVtWzOdTrHW5SJ08DV0HcHyLKijYofgsi197OG8GJIrQXpfJeWoZGNjkyObm4zH42QDpA0IldbC5/fOhz6PKITb0yyXA8bkLTYrksU6JZPVbgawXGwyfi/ytCgu6pmIXafXdb6C0Hd+yXA1hBw8KDIpgrBEhpDI/L7FXPwbF5hV9d7W1Wufs644f1hivt5uqLjcVNWvD9fFO1rnHy90OjzIIFBIVMwfaGRUiO5zSGRIx8mO4JLYlsvPNgsdW7KzzqnAOeK9/38Wjh2IBaW/zzRZQPchpjmrbR1tXSf42Tps3VK3LXPrmFu3307m7/W1+1+VGX7yjbCOr8si9Dd+7+Phr37/O28qpapyUCJ94t7rEJPtv3NonY5CISbfptl0ipDZoywXIrEUAho7c0ERs31MpA/+XTK07LylUpKqwusUTpWKiO6LV5cnRExML51TQ7vipJYovFKpfuNSSvVFpvv/5QK4XIS6ZFClxVJOSrbAzzOkdAKMeZPNuoj8/0pqSm0oBwOGmVTQNC1VVdE0ze1FKMORLAkGY0h5Q3TGpT70c5XknZX0R6PhiLXNdTbXNhmtjhkWA5CCICSExHjqNoS+yJHmPGmTFwfs+5ft3FK+nkSRnL0TVJlC8OhgR7Ggnvd/L6SfKQaf58oBH0SG3dKHywUnxDR7SgUo/Vm/+ZAKlYuCNkRa52lDQEtN0zTszGu2t7ZftpV/X1DsHJaXr+/6p1+86P6TN93zNLX9WEO8d3VQjjsLJqLswoFyoJ0k3wEIqXtLH4FOwYhdtQhiWRTW2y2RHdpDTCsaXCRElx1A0j0dsjdH7KTZIvTYdgyOEFKgoneepm5omxbX2lSUWkft3GS2P/kAdfxZXQx//2effrY9LELfxJeP7Djnp1IpjEz069ZFCiV7qGY0HuCDZz6rkkdTVTGSss+DcS5xmhIDK29ESvS06QC5ECUopisey4XIe58Hoak4dO7JKqeAClTWIqS5j15K7VwuQmqp6HQfy27Ny79fLkZpXpQfhNgN4WW/+cZ+jrPAuompgzDa4IqSQegs5m2e6bgeWlx+ncs0ZUFiC4YY+m5i0QkuaNal0ozGIzbWN1jbWGdQDBFagNLErrPw8UAn2cFgXXvSebwtd5ydOUI39xPZPVtLRVEU+KAJBmLUKCnQKs2+iPQQWoyiJzN0fUzmMuCzVsiTTFRdIFHQw1IxCh6PAKEICloUtYtMGktUFi1dsHUz3dvdu3L95cu/KfXoo//g05+3h+Xl678i8lpb2Y+aQn1v8OG+oPJcUKQIe6RK+iGVaf1SEmXK44pC9cSX7kk+KDbN692Jo/OaBu/Sve19T+tO97kgCt0XpmSt4rNEIEkp2rbFh0DbJkse2zic87R1u+ub5sOiDn9fFcMP/S/PPNe8UdbwdVuEXJQ3Z1W9tXZkMxoVhdaJ3SK8I0adpzQFo1E6oYeqxtl0Kumw4N7eP+20+BhQISCETKp9KZYs+UOChjoxYo7ZFt1QnKTV6YCjxVwmFRhiIkXIJXKClItIApXnOR2jTS4pt5fhuztZ0Is+6C1vsktsutQpZAiC9POkab9C6YKSdNoPCGwIWBcIoaJtW1prczHLw+AOliLHIHf+e3GhnUBIlNaMhmOGo1FPQBiORhRliRIaj8dlfpjPOUphWeez9MN0HgguQ3+JMr8M1yUKvhJZM5IdEWLI8xjtMVoBqRj1ptpLjtnpIOz77quDEBNrMCaIxfk0FwqZyZjvn+gDPkgisvatu7q3vbunXZi78bzeWBk3s529a7PrW08pWb43CHk4D/oDXv/ki+fb//0j5z47DOLLLsb7goAgIl4EZNb3IRM8FiQIEfosKqEy/CY7InY6sInsYBFEgmQDAY8nxGQjZTuhaSaVxC5+gWxgGiWRVHxkDqqLLrNKg6eaN1gfaEOkbh2xbV5Z1/r3gpf/2Bfmwz/zzBeaN9Iavm6LkNLFFV+1X9Bav12IuC6ix5hcBEQgCt13B9aWCSoKSUyGlOm0zYKS221JPsQUGS06FFj2J/FldlxXKHT2rlKFWcBv2Z8tdQP6AHQWpewTH2W3KaZBFyYz3pYLzG04+Z3oo12R7AumWPxMWScT4pI4s5uySIHShuFIIjMRQUmDMRPmsxlN2+JdYvmQqeRZioOMMkOBGqNT91EWJaZIM61BOaAcDDFGL2BMmVJliRIXF4VSLCk3utrQrU3Ic6XGp42BSK9HItOltdYU2qBUKoLS500lbwohJOdlrbsk1dgLldPhImbSQSBGj8vJl13BaZyntRbXZ8JkGr33iKRpmvrZ7GN+3vzTKDi/vV9X88L4bWNsCGLLB7Hz88+dnx2WlH/bIbC5pKN6DuI7oxDrQQSEikgdsw1TWrcoBELpnr6dNGgZehc5JbhrgbJCLGblT4pUsLRZBG6tTWLTJR0cSHzwmTabP+dS5xS9xxPxzlO7SOM8zseJ9P5zhfO/sTd373VCPfczz3yxeaMt3+u4CJn9ZjZ9Nga/i1HrMoKOEq8UCIX26UaNOg3enfO0LosaMylOZMV/NyOKeaP1JNquIqaOSKQNXC7Nh5KeoHNMlj1jTQp9oAhJZZYYb7KPilZqiSWXJux9V3ar2eLX9LvsRDbhFlisz/nJhDOR9RWIzBoTEBQSx0BJjC4pByNWVteo6pq2bXq7kWSKkOCxBA8mEgQymZoqpSkKk1Jj+/lVTjLtM3q6KVtiJoaQjEq7NeiV7SHkeIjUhQghCC75bzW2pW2aZGopVe/11Re7bO0SMnEpZCeHGCPO59C7HP3MkhGm94nZBKnrsc5jfcT6iHepGLnM/uuZeFGilMHP5+fdXvN3R6PxB//Zixcmh1XjD/cKyIm1PG88e86HdYJDRo+KHolGyoiSKQ7EKIlSEqkWTuayP+OEHPOeo0J8RESf9K8iEmUSMMfg8L7FucTwtM7hrMVnJ/bOjLQj+sQArfVYH7ABnJARz0Xt/fu89f98inj65z79la036vq9bovQX/vt99Y/+SPf+6yMckeb4h4ZFD76RMfOjLSYB5aJhlwQhaC1C+3NgX2827iFAJ9R5CBQIoAXRJUFapmeHENIwtRuRhUSlJf2ZXkAMlsUkpBNp+QiUEvIdHq/pQDd6vj71a6MjKWimjfJsLRZ9lTT7tcstkQohCTPrzSqEJhBSTkcMnbZ9de5/j0LsSNVpALTJYh2fEApDlrly9z1sQS3yWX7nHhrhDJ9R9qvh0ydj7PZDiV3Lc550IKiYxIuzdVS8Vep64mL9QkxOTJIlUXKMSRnihASBJM7J2cdbZ6P2RCwIaTuqINn8hnaBo8PWOX5jB6ufPafvXj+sAD9EVz/2/Nfnv/lxx96aSDUThTqnJIKkZ0KJIkaL6TIRAOLQKNloiOo7j7o5pv5GZA5HkR0z4VWSJFSfIVIB6Hg0n3W1DW2rmmdI2QqdpInxOSpGCUharyU2Cida5ov1luTfzQcjn5Vl+Yrv/C5F9/QurDXdZ5QUQ6vYv2rQuknIyFtRCFk5kzWnXTiTmNwMSKcz51Q52CQx9RC9Juf8IklFzJu3KWHdgan6fPZ5yzP+2XIN73sIJ+FQ8Ji+pC22UV42iKTZ5kKflujE+Mdu6FFouki1fG1beVjdqZeUFQTKw2UMYuIYiJSaTSSqARKB4ROUBRhQVXv9H4hbwJKqhw4x+LfJiaftmyv0jkciNjZreRgvOjya4vZTikcfN1Zk5MGvom9J6VmODQMBgMKY9BS9+/7gYCznouRTERjiJnQlH7ekAuRCyHPd0iMuBD77i90jDpB76TtsqYkRDkptH7Rx0PW2x/lNW9DtRb1XEtNCPkjKiIqb3OKGBRCGZQqQJrkvB4EQsncMclFGmrM4YYxfU2QAqLGKEErPTHWOA+tjbRtoHUkR3zn0gwp49JCKryXtEHQuMhsOjkvK/vPjCh++Z986eJLhyv3Oi9CMXLt2iuXPjdYLd9ltDqiJCmLPkq8zHMXJXuYRmcYKZKtXsICBpKZvixibrl7nYDqBa0HNti4wIrFYtrdfyzbvIeQPKvSyFzcoZDEO2ph4i3F5bWK0O1+V+GApsd7f2BW1HeCeU6UDEzDoq+SIg1gBQilMEKiOpNPOgiR7P5NTkIVWWexlOWTnSaAfrjbhYxJIUCmeZCIiuTKlQkFXfRBCMzrCuc9TdMym8/Z39vF+cCJk6c4euwoRuoMrcoeGl12nojLlkzdzx8jgjTP6SMbutfeOWULkQpNWDLAzO9vNyeQhaadN3vBhS/+4vPnp4fbzR/N9SfueWhlez49vdJurKuoaKWm0CVGD3AyFR8VNUVR4pQmRIERmqhM6sSVImT1qtKd/VS23pIepAFZQO6iZBRIC8SK6AUtjpm1WB8QqqB1Dus9UUiQmnndsrM/Y3dvtj/fmr3/1JEj//rj29cPC9AboQj9d7/yW5O/+UPf+T4Vwo8bPTjSxAYpIyHKniIsujmAUkgfMDoVIeGzt5Sg3zwPwluJGRWETESFW07mt6ZwiqVuKRWlzLKLmejdsaluzXrubD86D7qlwthDWEvMuOXi0/3amSgmG51sJ+N9nrtkUW33PeNibpS1lQfKopQSguy7nARdJJYfcjFL6/7dxKvLpPDcIZE7jeh9+o0Pfdxx9KGPOQdPXdeL3JVcPBvrkrbCO9rgqOYVddOkv4dgNBpz7NgxTp8+jQhko9Qklu16T5mLfhc/0ZNQ8owsrXNY8gQUWe8Te4ZcF9HgQ8BF3xuldl/jnGM+n+4aVxyy3v4IrnecfXAgQji6XVdPFoX8i96UZ9qo2G0jlfDIapYCEMmHJVMkAbTRDIdjRqMRpihQmr4Tl4vWOLsj+LTODkJQNBbqqLBmiMPgg6JuPFVtsUHgbcR7w7z17Ez22NqbsjcPtM5jXYglXFhx8eXD1XuDFCGAYrRyqZD6ctO6B6VSMkoPMXU9LndDSU8DSnq0kqmVFp2NTehpv0LmLUxKXFbQO+GQaJz3dFpPGULyO1vSxWgdDxSh5da/U14LsYijFqLrBmS/USY9T1jk3Gf7Gr+kV7gTNBecI3qSf5vPnlXdbEjEvgAuOyf00J8/CAF2VGshOjp3ZgkuWQ/73Dl2sKLsCmQ2jZRSJmjLWbxNjgq2adNcJ3i886lw2BYXwYW0ZoEURli1DXVjmbd1cgkvDIOVDZRS2LbFKMWoTHEdRqfY86qqqG3KL0onXZFD7GQ2Ngh9ZEb3HsRMiuhgwO5w4ftspMTMcyHgnb9Fw0TqGGO4GaS8ebjV/OFejx0/t7E7nb69xf5QiPY9q3L40JdfvbIeo0MoRYhpjicgO2/o5FrfOY8UBUp2gYwS1YnH6Zx8U6hkLx7LrvVCCJxPDiBCKoL31E2Sdwgh8NbjQ6T1kZnXtLIkFI6gJGgXfRNXGyEOtWBvpCLkhb584aVXP3jqwXsfFTGcVFItOhhlUAGES4wXrVXygYtQKIET4MTS/IJE8e6EqcnGRaZwLLeY32gF1ocUKy0EQoILLg1Y8lwk+s5zLb0eIbO+CNl3HoGk1hdRZAfg7qgesp9VKgl+CQrrHKf9kmGodRbrHcEtNDZ9CLHK7uFS9q8hhpi6mBiTcaOIvb0QefNeMABFSp3tSQ0pJM6GbhYkU1HOXytjxDY1TVXR1C3RB9q2wbdtEvPlQiRE0iXVMc1gprNp6toCyKJk5hSrx88hTUGUiUDhXYOUFaPCMBoMMFEyNAXFikRLgZjPaQSJwBBjFusuoNWk66AX3WaRVrLXCSFF8WZvvC4byLmIFAonY2IJ5u9rPYSoKymKi1IWW4dbzR/e9fDRM4Obu9tvm9jq/xKMfFtZFMdsVZn9pk6QWhaF11X6fVGUC3NgITBa90SEZV1fOjApOjvBzixQ3AaBp+PYcgx4j4K4TqCd54NmQCE9MgSctYMY2jNB6zVg93Al3yBF6P/6S78++X//+R95H1H8WSHUSaVA+M5FIJEKZI50IESUlAQR0FKhlEB5sKl6LGC1/sQPKoCTERnSiVhFlTqBkByyQwg9zbj7WHZy7j8yzCZFFtjlrigQUZ2lzi1fH7Ljb7ilCLk8oG+aRKFug8dFj4gSLRXksLhASB5aUi2SJWPoTT5VFAip+5TJFHucvocSqndkaL1PkIck6ZxI8ckCgQipkAHgPI21tHVNVdU5Uyjlqnjn+1lVjGCdZd627NuAGgyxJPFsUQwYbRxB20CxtkHUBhcDBAd1RWgsK2vrrAxGCO9QRJTWuKKgdI6IoMX27/cimGxhFivzASAszXniUtLqQfcGj4sC77N3XmetHiUEuSei/mKUsjrcav7wrqppjk1t9eNO8Xal9akoBE4oQtbkheyP6GTnMG9SCGNmZ4ao0sFxCXqTMQvEI7dMZcWB/086oIOfX2gEEyGls/IidqGO4D2EKIqIOBqFGByu4huoCAHoYnhBRS4Hwltk9nADMvQjMEpBVEQberKCymQFmYN2ujjgHnXK1GMf0qYdhMCHHNUcBFHIA6wzsSRqS1TvxYwnQW8KsudY52NGDMheMCuWClDsZyTdVMP7Lj4iwRBN09C0Dc77HDshsyBPoiCrPrvo6mxsL7vOLXkOq9z9hEXflDomIlIEoktRCkOletgxdLAF3Twow4oxUjvPfDZnPptTtw02F4WIpImOurY5rlvgo6BGUUvJuCwZDMYMhkNW1jYZrq7SonAImpCIE001xbsW21asjE4xHI36067KGq3BoMxar0CwB81kl4ZwSwQKbj8sdAeAjrwhYrYzCvmeitnOReKa5mawPPsbz3/psAj9IV5N2560+CelLo529GqRafcHotMz1LrsvbgMKd9aYKCzbHrtK9z611hEv8ecSdRHPeRnNzlrpGdTxKhCiIeL+EYrQjb4nd3r159bPb7+LaEwx7qWXWuNcw3epVmFEqkgxZhYMsZrrAuZJpxuNMmSQFSQ3JJdTEmoQWJDQAVJkOkEFIREOJ9w6luKUJoLdeabWafQ5QwHcnZRJ9A86MLdbY5J8Z+goLpLLLU2e1SlgDqhTSYYSAiWqCIKlZhpnZebWtCXVUclCImAUZYFiICmO/FBdDkryMfeWsiYEi1zWqwQOO+p2xrbWBprqeqKeVVT1y3WO6LUtN4RkVTOM2tahDKMxyusrq1yfHWd8coqpihp2xahNdoUNDZ5+oTGIqyjUAKhJd4o1jY22NxYYzQcIGXu7rJrggkG5yOtdwh3e25czELYA9opDhai5TXsLP1FTrztXMOz+0Tt6+bLEfni4Tbzh3edXT0qZ/P5RoQNKZXpZpd3+ljEphxkRC7HoHTX8u+/mvbuVt3a8v/HvD8cYJh2M9B0/4SIqH0IhzOhN1oR+j//41+Z/p0//yd/Z/342g8IJY8lFbNH62RomTzF0rhGhWRmWRiFDwbnHJUSJCZCzrDJJAKRM6JjFEjvUCi8SnoB7xM85WUSsXadUJ8FLrNsv9MfdV50OZtRiIPqobicY7OMOYdI3bTUTUNTtwnusi22bVPRlBJlHSiBVgVCqVRIdRKPChERQmZRn8oiPZWhQUmIjpvXrxKjh94FO9GZE4FC9nZFnbi20+DEGGmCpWksVdMkn7UQmdUVs6qm8Z5yvML6+hGOnDzDXaurjFbX0EWBVJpyNEyxywSUbRFK4qNEtW1ywNY1xjraakaYOYieE8c2KYzEhYaIYCCGPSVcKY3W4cCGc1D8G2/5XOite2Kv/wlLVi1dtLdHkrVE2SEda3cU4qmo9CEp4Q9zxhuiCDGUCFG+VlG4tWjcqTjdqfAsf7zWFW+RV9x6Dy0zVnsmbHdwDcEH4pRIe7iSb7AilHBg+Ww7nX7BGHOvVno1RI+UySk6dKamEYgOT0RJhTFQOkepNNa1maBwS3HIyJbLWUPSSmSnb5ESKyKagMz2Ml64LCsSOEe2k08miqLLqQnJm+42H7goevZVIDH2mtZRNw11XdG0yUKntWke1CW7FkZjTGIHKW3QUqIkKJEKq1GC4C1tU9G0LbZxtM4nO5rQont2W9YYxWyDv+xCnGO2ISWOtk1D4zyNs0xmcxrnMEXJ+sYmm6fOcvf6BsPVdYrhEGkMxgzRwwG6KHFEnE/hgh14YoLDx0jV1AwGA2KIWNciHLRtTbQ1AwTHN9YZlAatJUarTIFXB07A4pb3ltvmPjEntS40SX3xX+qGrE2zJe9dhuJCFuca2vn+JdfwSTEs9w+3mT/M5zhGH7t8Y75qAVo28/1anc1yIfp6v/5O/95X+1ohhBdCTInxsBN6Ixah1vmta69e/zdrknesbx5f7QQwWkti0Eg8UmSqdgSlIgbwhcEUCmkFNsQ+OlF02SEdnTkGbBAI7xA2O8kHgQwSLwQyU5290IkUkWLjsr0M2VYkCyaD7Pf2zqU7QXiSbgoUAliXrOHb1tLaNAtyPsUstG2L9x4pQBPS91GK4NoUP+BEThN1tLYh9my6DCPGLqwtZlIDfXR2BILwaYYVI60LtMExnddpE9Yp8G68vsrq6gqrUqGKgtFohdXVVQajMboYIKRGmQIhNVKn9FekoZAphM/nH3Qy22dvOmd/OuXSlVcJ3jHZ3We+swW2ZSgkJ9fHHD92lJGWqOAJ3maKdOzdt5fbyjvDKcsFv6Nkp8LiY+gzhELORorBYX0iVkils80/BNduV5PZR1Sx9ty//MILhwOAP8Tr+nwnjDAuuTZ+41y32mjF2wTiEcBLIaoIh0XojViE/m+/+q+bv/mnv+cT4ubuF0Zrx84qKYYqAl32jlREFfEqELzEC5nSu8XCCbsLr1ocbTKTqgseEeCiRIaI8hGv06dlFPiQjHuX23YhAkrl33ufBuki61dEB9Utt/6Lv+sDySnAtn2KZ+d+4LLPWQSkUCnvxrZEBHVr6Uin0QdCcDjbpCLXDeSFwMcMs8XkEuEzPZqsgZJaI5RCmAIzHDAoC8xmRBclyhh8iKysrzFaX0OpgmIwwBiN0QVFWWKKElCpm1LJXbyqKrZ3tpjN6t5+x/mWK9eusbO3Q93WXLl2Ba0E9f4+oq1ZNyV3HT3C5umj3HX8CIWQyBhQostTSuLXuOwYxO1WR/EWjVWfLZPnRLfOhLpTdvIIC0SZCpVDEpvmZvTio0KqQyjuj2LDh4aFhcdtPox/kA5mWeT9dfkwvgb8d4eu5w6dWAwCUS2UeIfXG6oIAXhhLrZz/ztNUz1aDoYPEWNv1xNcR9UGpQUqe4lpJSi0QuVMBankgsVGwMaIVDKHnwVEdEgiToJTnY9aREqT0jUDPeyWBT2JoZY1NComQkLMR3ORzUSz/BMkOB9pmhQJHDOPLUSHz2FrnQ2R0TqJ6VqHVApbV1hniUItYdf5O/dO1SKHtoX8nimstQipaFubiqKSDHSBFJphMaQ8epT1I5uUwyFmOESbItGmpaIcDHPeUJexZJLLgIsombq3GKCpa3Z2tjl//iJXr17DWsvly5ex1nLpymXmdY0yktZaZISBgKGIbJ44wqmjm5w9eoSBFKho0Z35aIgpMybDnwmaizl+XfZODB3jcLkLIibm34Fo9q4jynOhpml61/CqrtHlkLZqrVHyRV2Onv/tL58/xP7/CC4hRBMj/tZO407d7fJ1awZXd2hbnmHemsX1tTqeO33+1n+7mw8RCULIZsnT9/B6oxWhv/Lr/2b2N/7sD/7O9VevvvPuh+8/EQLrBI8g9gF0IcoERSXJNCEEdA6Sw/qFpidZRi+crrsANyI+JrGmdgEh0kaXRHAerxTS+wMnt25DTJ8MvWNCH8fdCVCzUt86l1wE8jwKLVFBM5QSpTRtPacsS5RSXLl8hcvXrjOZ1AxWxgiTyQlK5RgJSQxhSSKbCp7UCq0LRGFYP3kKrQuKInUxZVkwGI1SJLlKAXi6LPARoimQwyFFpsoCWOuSJ1+Eq5evcuHCRa5du8bu9g7z2YzpdMrVy1eYzueJmSgEw7KkquuF6at3OA8rQ0NbWQZK8OaH7+XR++7l3pMnWBuWqOARAWRUmXTBATguxOR67LOI99Y50DIxgazt6pwRXH7PnXM4m/6+1ppZNUdIhTKa6axGKrUlonxGl8NDq54/ujLUZjz7Nc17v1ons5wIvPwcfj3f59bO6avBcHeqYULQRsFhJ/RGLUIALoqLTJpfrmfVWwbD8q1KpE0vSgXeo03SrcQcDyxixDtHWVTopk3ssE67k0/a5FOy7ELt8HgRaXLXrTwoBDEayGwynfGEKBJNWkvRQ3qyNwkVvQdCFCk+2tqUZeNCKnYRkTVLMXc2afPfWF/n6OYGCMHurOHKzgwhDOtrR6EwKFOiTIHRydJEC3pdlFSGYlgyKMeooUEVOhXjPvdIoIoiW9QHTFEwHI/RpiCEwP5kn4uvvMqly1eY7U+Y7O8zm82pqoorV6+wtz9Jcdp5oy8KTbCOUim0Nklk29YMjULHZLMyKjRNUxFry7Gh4tEH7uGdT76V00fWWDUaGQPetUhZ0EUU9VqfTNPuTFK9D7exmWJnRtrlLC199Nb8XW5Q8LjgsW1DjIG2dtgoCNpQCnlhNrfv/40vXdg93F7+yC6bljXeEQZbdos/YDm17P94h6LztbqgPwg8d6cOKr9gfwjHvcGL0P/j1/5V+9f/9A88fenF8x+466Fzd0utjsQ+RP7/z96fBlmSndeB4LmLu78lIjJyi8h9rcrMWlAogSBIQigSACkuIgmKa5MUJVFDaVrqFtXT3SOazWIaa+uesbYZs7E2m56x0chkalNLpMRNItVUixQoUQRJAEQVyULtuVRl5Z6xL29z97vMj+ufx3033d97kZmVlVl4DgtkVkTkW/y5f8v5zncOK2ytOSQcLMZsjCQxaCVNdPsZBpkqzKpQWmXTxWjg1AG0NYUwqkXGDKQBONfFhcpLxWqS/mDFcqpD6DiYNWCGFww0Jx1DWliZUgUVGGUnBtqF4BxJkqDVbGB2po25uTkcOXQId1e3cX1pDRvbHcRzexE1ZqCYhFFAxDgiztCIYjQbDTApIaQEiyKoOILlEkxGMDBgcYJ2u+3gOcbR7/SwsrpSwGYK6+sbWF1dxebmJra3t536trZQmfPeiaIIyijEACScTJA2ALe20O9yS7ARB4TgaEQC3BikvT6SRoxmHCGSAheeOouPP/M0FvfMIYGFNRmUNogiWSRKCcMcVZ6LQtG7YLGpgrxBycf/0xiz0+UWmn4wGraQYlFFAiNiglYWXMSO7GEZhLWrWXfwhxDx69PQ8sEi60B1N1HX1VQlpaqkU/f33XZbVc8NcjfBtBP6hk5CAPD3f/N37vw3f/Hbf0MPBp/Jmo29Qhsn6EF6YiRqCAEOC2MiNJLYOXXavPCuL+i7lkNrWzih7iw50vyAGwPDOHJV7AwoU3jak32ro0kbayA4c06OZDHNnIii5Q4eUkpDa1qiLIy4LAPnQJwIp21mLZI4QbPRQBJF2L9vL44eOYzVrW28dfk9DPoDiPass2goYD4uImgZO6hQShgpweIYvBGDC47+IMXG1gbW1tagshzLS0swWmNtZRWd7W2kaVpCimmaIssyqNwlZwEGWfgyaZVBcmd17pwnLZIocuddMMSx67R4FENwDpWlSKREu2VhjUar2cKFs2fw3DPnsG+ujVYsYFQfHICIGGQswCIBI5wG3458iiNWONtv5cRGgy7o3j0hA1OKkhbMQWWgtUFGcB4sVJYBnCGOYqyvbdw1HfXv49bctAv6YGdCCvZehpkf/KvUMCbZAarrhCbZR/LV8sPl2PIxreXTT3CahFxwFNFb+UbnjxIZHTKcHZWCOyfEAsvhXJTLqTIyaCYNxFygb3ZIA05+ykFlplCONgVDyllGOFYcuEtGSnMwrsEVB6wqnEfdbEdI4QzkbCE3wgBbSPsww2CshjJmSDbEr/qkEDDWItcZpGig2WghacRgnOHgvj04e/I4lldXoXWKLB84ooB0Uie0PGsZQ641tM7RS3swm461t7Wxge1uF+trK9DGYH15BVmaYnV1DUoZJBF3VHPviDggOXeMOmsRMydyKriA5K7xjOMIUSEDJIRTaDCD1Nmfx7FjJeYDtBoJZhpN7N0zj5OHFjETS7BsACYTRAyIBAeXHBAcyhpwvSOeSkKzbq9HuZ0etgPXDQehYF8ILgEZS1YSrnMj8oYquidtLYyyW20u/jhLotd+88139DS0fKBpSKOC5lzV/dTAYg+0DzRJAqr6GWOMFUg8m36G0yQEY+zS9lr3X7Va8XO55PsQN5quu/A2q4vhNhCh1XbaZdvd7s64gMzovL0SxgpHzkLfjdx0clYwsLTzyRFggMpL/xppLLgAtODgpuiAUOwPcY8uXMJww2Z6jDFEcYSkEaPdbCGOI/c+VY7ZVozjhw6gc+EM3ru9jH7eh7IGieDI0g44ayJDDjWwSNMBut0Otrc72O5sot9NsXz7TmFpXQiVMpdgIgYkkSiSNnMwHkcJf1ljILkFh2MgWgCy8F9CIhAVrDzJGIQ2YBaIk6bzdNIGTGi0ZuexcHAvTh49iQPzc5hrtdBuJhDMQiCHtgqWyaIrVWA2KiBMAcsYaFVVa40sS4eS5T3EBOqOjBkyJdz5sp5agpsdiThClufIe/3bsea/H0XRVDH7g05BgAKgLZlx1SSacAbkkxJCOZ8ycVBBVp9x7gHTrLWlIREzqOyEitfCrbUJMO2GpkkIwN//rX9v/q/f/51/srnc/RdiT9IyEB/nQjRjWEjGCpZa4TdjBVoNhnYjxnYk0Fd6R1+sUAmwpvg31ilIG8YK7TgDGAkFekyDjGmIIhZaMAhroAyHMAbCFDp0xc4QM8XNI7ybBBhyYZVCwjifBgixY1McyRhy1tlaRzICf+osMmVwe6ODvs4h8wz9NMPd5WUMBgNsrq9jdXUV291BsUrr7vCYOV29mSiChUEcxVBaF0QGS0kdQrouUmsNcAYmnF+LY/5pCMYcHMc4YinBjFMfbzUSCMthVI5GHDmKtQTm9jRx6vQJHDy4Fwf2zLvZEVxiMzpFqhRkVDi8MgnBpBOvLNxajbFQRsEIAZXnTg2iMNBThahkOA8q5Xi0dnbhBsi13fEP0jm0JjiOIRuk4FxsRMb+kbHiy7/2xju9aVj5wPE4DZeIbJXixbhOqLR2x2SqCrvpkixs7VwJDNxa27JTSG6ahOj4P/3W7278N9/72V9NBqlpL7L/rYyjjyNisbGq2BeKCs8fCwGLRiQQCY6Bytz2vGUQXDhWFYBICjCjAeYM4yxnMIJBW40IwhEWjHa+PrYoqhQgIBExXsj1aAjhLLlJGofBwio3r3IqCkTatkUn5qSAnEEfh5ACcdyAMaTlFoPbFM2kgRcvnMP8jSVcv3sXy+uruHXrFm7eWsUAKNIpIHmhmC0FpBCQxknoFJrE4MyimUSOiUc7NZIVIy4Dy3ZckSxnQCRpTwKSAYmMEHMOKTgSGSGRAk0Zo91suGTJgD2zbew/sB979804RXNoCOEWZ9OsB84BGUtEUexmaYW7KzOF4oU14AbgUiLPdmSMlMqKHa3CIFDv0O6tMW5fyjrYUxkLpZwmnDYGKs9gVO7eY7ErlhsOkedXhBb/GiK+Og0pjyIHwTAgt9baKlHSKg24sCuhZOQnonKPyI6H44YSnN35sjXzJ845NJjQRs9aa8T0U5wmofL4v/zb31v7P/+Fb/+N7ru32s19zUY+1zrfbkZxbDmUyQuWFdAfaPSzHP1c2TRXKZeJZhaNQZYKMFnY3THEnJWuohq2UJlmEMwAloNFptCAY9CKgYM05TymDmmcGQtmdQELsh2fLQxf/w5BoFkSwQ6sNKiT0lkbR5lCxDgOH9iL+dk21rZ62NtuYWt1G7HSyK1BbtzcI5LC7TZpg4hxSAZEvEhqZDVhnEupLGBLzuC6keJ18ALWsMx5sAjG0YwitJoNtBsNNKIIkZBoxBGSKEIjlmg1mmi1GohiZ8MsmTOk48KRE/IsLWZoEeI4Lve0nPFEEQAsAFvsUWmNLM+QqbxQuh5WPgir6CGVbLjPMC9EYVWuCtXyomtiAtzqO731rd9qtfZ9+ddee3swDSmPAo5jtvCbtKO6nrAT8YkH90vDDuc/4XMQChF2XsYYcMGj3Jp9xhg5/RSnSWjo+O/+3e8v/72XPvXL+e21iBvzn3A2e7ov+B4hYgnOkRlgdW1jbXVlaynvqZtC2TtZv29TY04jTs5HiTwgrOtOXHBybqTQzktHMAldrAgYQ3RuJ6JtDAMzZmdZlao1ENrNd6R7KAFV3kDFAL4wziN7cFWoOidJjN6g76wZJEcUtSCkhFYZvu0Tz2JtfRN3Vlax1eki004ZGsrNuKLIUaq5tZCcQUqOWEaIZQTO3WxMcGd2594vB+MMggFSSgheuLUyjiSSaDUaaDeaSGIJKQSiSCAREkJyNJsNNJoxCh0iSCncX70FU7LhEMUyLDlmlsGlSPjGWhitkKUZsixz9ujgpe2Cn4RMYRKoqBPSjgiS5ylUnsMq2h8qnDYYh1JGRcBrrDH7u4zLpemd9Mg6IUuqA3V07FHQWRWDbVwCC3/Xh/H85/OTkP8crjDjMThbsNa0p5/iNAndc/w/vvTHt//eS5/8n/vr/ZvM4PNGsBMiSuYs47o3SNe2VjbfTDf7X8oH+qa1fJNZIFLmBGD+emb6350kjcPMGigwCG4B65xajXZ0bF5QFEpYwDoFN150Pj6EYDyX1ULVDKb8b/9GgKOZMTcXsXDW1Uq5fRgTucVNU1DIIykROZk2WJOjHXOcWNyP44cP4ebN27h28xa2trvodPvY3OqgN+gVauAWURQjlhGkFIgjgUhETjWcM8SRgOQCsYjcro5wrqvOn0kWpnYoZ1ONJEazEUPK4veEexwpOGQUFcumDDISsMwgUxlUlhUJMUKcxIiiqExInHOnOk7ae0W2ttog146arZS+RzHbzY3M8M5QURA4g0Bd2jXQoZSFthzKAjDqJsvx2yJqvfHLr701lWJ5ZEnI9brFn7tiulV1TFULr1UwXlUiG/e8gYUE40IeBOwBAO9OP8lpEqpIRC/f/YXPfutvZBv57wvBFoW0s8oi76X5Zj9lK1ok6//07YulHthPP/v0tSzP1hOgk2Pwl2Qkj7rBiFMDgBWFta+GiAUA47olZ/3sZinFxtE9F7513qTc2aCWjDNwpz0H5hKZ8+HeucEs3D5RphUirRDxogrjEkkcQTVimH4PWdoHY24Wo6FwfHEvji8cAOMSW9tdXL9xE7dv30Gv10OUxI4uXjhCCiGRxDGSYq9HcNcZNaMEccMlKtcVcURcQjDh1qEYwLkAlwxSCLdIagwgWOGMWbABhXOxNUxDZTmcB5gtjPMixHFUdkFDN3wJUVooo2EsMEidx5LWbk5nqpxSAxhOFSQER0TQpcqCUgVDztlVbCBTX9Q2+be/8vpbU0bcI4Xj3GVorWWjkskkCcKHzKo6n0lUFPzCserfU3ckhEAUR/NMm9NPHVh45fLK0pTKP01C9x7/99/7Sg9AD8DNcb/7i29e0gC+/uPnz/y/pNGZYvZH40Se0IX3DQQHZwLcumBr4XZxrHXq2I6oUMB2XN+ThPyLvxRZNK4zgnXU7SGJEpAmqkY6GLgupNFw+zJ0E0QxojwFrEWeD6BMH0nSQEM6PyWtM+xpRph76jSef+osjLW4u3LXWYb3+0gHqZPakc7iIpJR8SUQy7jogkoKAzgXrpsquhPGC8iCFUwiKSAbbrajiWARSajcIM0HMEo5AkPi7CGE5PfQbUv4EgCMO68GFplSSAdpYVGhyyRUJhivA9LGeDbMbjk10zlylRZ6cwZao3ADFGgy+3puk39mefTO9K555EfEgIRxzv37o+6ogufGqW2PMrir2gfy3FPveT1DcJ2Ue6zJXjTG/DaAjelHOU1CD+X4lXfefedHz535H3Wnv5la+1dFHJ+BziHgKnsGC6MtYDk4eRAxW9A5OQANxtQwxVQMs378BUpKUHQj0KwE3DmjamWQDjJEMi3N7DicgnUcayiVYKbVQpZlyAcDpIMuBBOQPIIUzgAP1j1ODoOFffsKMVDXjQlWOLYyN3AdpKkzygPfsaEoqKokHFomUiHApZsZFVM0WOE086xxSSJPM6RKwSiFqBBSjWMJIXZcWylAaBoOF9bj1lAnpJArR8vWnkI2GdPRlyqSkSG2m3L0baUNlMqL5V2nVGEMh+YM+SC7mzDxu4zHX//lr39dTe+AR3tYa1oMrCWEEKFMT9XsZlQSqUsyo7qgSWndVa6uQkYzVulPKq0XpklomoQe6vFrF99990cunP3HWW8AMPuzMo5PMRgwrdxMh0ln3M2cpYBl1iUpMEBqCG2GWnvDNDgP2nwGALyE40Kr4XLhEk65epBliPIIPG645AJAG6f+HCcxOLOwRkH3cwzSHqx18jORbIBzCQiOGAxWSrj9n4J4YeFgxMJ9NIlkYYPEyoRQ3nhCAGKnU+GMA9wWqgXFsi+zjgjBAG2cM6yyGnEk3esRElLuaOkRg9B4ZnSueWSl0Z7KFbLcCb06m25begaFenHG2w9yXVExE7IW2unvOzUKA+Rap7rb+1oq27/1y2++MYXhPoTDGL0XDHPDQ/9qQdKqhdWHCg3WWDr4h2/1LaXkuRRP97uDT57dv3D9yupSf5qEpsdDO3797SvX/tL5M/+E5Tm01T9jI/GUtRqxjApmFsCZheEALxhshjHYnIEzDQ6fZcNgLAczhZcqM2BWwjDmfs9YWI+JY4yzgOCMwTKL3FjwPEc0yMAhgAgFay2CiCJEJoaxGrFNXKVv3U5MP03R6Q0QRQmazRZkAdM5Az4OKwQE4ehDZPGCOOtuxcJDCADnsLxYKLe2cIx19CZrHPsOTEOrHFlhkcA5RzNy8FskJKRwhIxqhWRW7OyQwSCQK4VBmiFXurDAcInJBiQEX/1Aqx11bE17QdrCKLcvpMGhOWAG+XWu8RsZs29Mr/hHfxye2y87vc4JMDbjQ1/OwNAOwWBVHRElg3BHaJymXEjTDh+3xkn1ntkQYww5Fwua40eyPP8agEvTJDQ9Hurxr955970ffebM/8TSQZ8x+3Oas6cypTiTDBwChrlERLMbBgYuOJRS7sYoynqmCriKOyM9xgRY4TVUVWnZwnLCWuOEVhmDynPnyVPs9iCOwYWEEBGEyMFFBM41Gq2WS4YD59JqjEaqU+iBY7QlUeyo1wUTzd3ArJxDsbJNYx6F3BmgO8lxWzIDLSvNY8GEhFJpSQSAtZDcLcjGUYQoikpb850dKNqZYmUXVGQ4JyyqLDKdO0UE7MjsWFMhw6NNoYpddD/F7ChXCnlhdW7BkCmLXFkAWM+2u78V8ebv/ut33v5AlBFOHjgiGSAZY8LtfjHDGVMXb1+bWkK7JDJrrP4mEcmZMHHUJaCH2e1MCsOFHRi9NmMMhJRNHUefzJX6rqcOLK5cXrm7Pk1C0+PhQnNvvfv+jz1z5pcSq/Mc9q8oxp+BQaNQ9oFgjidnii5AFLHaCktXbTnjQGQhmAQzzCPC2bLjsN52ty7EO1G4qyqlSs05WKDFGIQUhbU2LbpypANHTpBRjIYxyNIMgzRFf9CHynMkMgFjgJASURQhiWMnD8R4KR7EKRsV+0nWMrDCrsF1cUX3oY3rggqlapU7Vf6IC/A4cqw6SnRmZwfIdU+s/Hsp4cV40dkAmdLOc8loN1+y1i2X6jr4zZQdkTIaqiAk5Jr+bpBpA20FLDO9dGP7P3ItfkkBVx/0Gjm+9wizxjSs0TPG6LaxZtbCzA0GnXkwto8L1hJcMMFFXzCxdvbgkSsMuH15+dY3dMDSSu3V1nxciHimSpVgt/DZB3XUJUhy9Y0ajcO6P/ipTOWvnT909Mvv3Ln5DcuUmyahD+j41bfevf7jzz31i3rQu64i/XdtlLwYcT6bGwutDaTghV9RkU6YhYApF1Ppe2A76s5SynsgATdDGtKncq6w1gDFkL7T77p5BwyajQYkhzO0s06BzmrnT8TLRVcOGUkkjQR5nqO/3YfWBnmeIR0wpFFUJAoBxgSkFIU8EFmki7IT4oWSgrPVtt47dEkhjmSxK8RLskNZ9VoD7TshEwvOAtrQeXJ227kyhdmfKckHpjAJpJt/iI6t/USkyt2qXCmovOikLIMxHBbITaa+ynP+/zVcvvrbV9/dtR/Msb1HGkabttZqVuv8QKe7eYAxe8Yye84ynLbAfsb5LBeixThrMMa4YtZy6Jxbs6Wz/D3k+n89Mbf/t4UQ199b/8aj9x7dt8B6nc5ZLuUJLkQcDv0fZZKZNPnQjJeSEK0WMMZiJOaZfq//V0UubgO4Mk1C0+OhH7/yxuW7P/rs2X9rB/1lnff+PmftT4pIzimHUAEAlDYAAyS3O2wxFE6pO0ztGliAgXNHHfbnJcYYRwWnwG00+lnPLanCoBnHhfQOh+ASSdJ0r0XlDjOXABfMERgiiXbSKKRrcqjcGcJlKnWJwABSRoUpHS8SSuQgRDAIOBiPFUlLSl6IrJIGHivVq5X1MfuCz+22XGFLXS8yqXOdjrUGudbIc9fNGKD4vntMxnEPEUHrHTp2nufQhV9QplQJDSqtoa2EsQL97e037Xb2DxmL/+i3r783kTTPib1HmNa6pY2e11od63Q3Txvopy3MOQOc4EIcFFE0L6VscSEajPNECDG0/+QFV92znVNb3c757X7nwkzU/scn5vZfura1+g011DZKz2qYTzHB91Uxzx72ManlwziHVn92NeR5JKMDJlaftbBfPr94ZOWdu7c2p0loejx8aO7NK50fee6pr7Js8N/qTuf/yGbYNzEZ7bOkPWJd0NTWghleJCG9c9HyYuAf1N40l6kIWMGN4L60VcjyFJxZMGucUKi1EEwA3EByCct0KXvDAVju5G+s0UXHwmDjCNo4lp2xBrYw2WNFAnJDYgnBndWELPaIyhuQu3atZKwVBoCkAWkKHTwN96vkrcTsTgdlC0sFbQyMBjKtHIXamp1kVZybIfJBQcfe2QXSw+oIeue/jXVsQJWm75utwS8zJP/ht29c3R71WZ+cPyyV0e08z/dvdTZPDPLBUxbmE5axj/NIHJEymhUybkVSNqSUjM5XeTMWUkQUtKIoos9RpGk6ZzhvpVr/dJp3L7Ty/i8dae/5moziJS749tXVu9lH/V7K83xPrvNPiqgxNwnEVmXnMGnyqRI43S3M53dBVFzRn+V9HMVHM5X/MFf5nwH402kSmh4fyPHrb1we/MhzT/2Jzdn/zfYHf0tF+iXeahwBZ+DGwnAGawDOioXWQs+acwPGjZPatqayuqLsRDeM1tp1HcXvaK2dDYSxsFkKGLcgayKNJIogCtICZwySSxhosELpAUUCMCV8xguqsoHQNLNyAd8JRfCyu6JZDi8o2uCOLWeKXR1jC2KAdcul9F44ODgzhSipgSwDgC1p6dpYKOXESI12NGpbdElEaTdwSV4X1tw2SEbuS5VJx9l+e12SZYAyt7K17r+2ufjNFLpSG+7k7KGmMmomV/mh9c2106nNXlCwz2vgaSn5/lgme2Qcz0RRJGlATcknipzyA32m1AXleT5kG+8VGVJKuWC0fikX/JmOHrwjTfZyIuI/OD637zIXYpUJvn515e5H0j5a6/yIZewU47wZFl8PqxPyWW1Vf69DJUKW3bgESNcBY6yltHoxzfPveOrgoeuXl++sTJPQ9PigEtHWjz3/9B+rPN0QSl82ef5jhouzEYOUVgLGwPKCNWedmI8GQ8QYIlGwwKCKCx7g3JZSIGQVWu7nAA7C0sXuDNzfDaOE5jTmtNGIuITkDJBO682t69hCDNUlBRFxF8S560AY57CFc6xjwLGd5oPxYgHXEQmUowEC2u50MbaQ0LG6UI8wzl4BBgy8yFcCnFmnLm6Hdd/crEbDGudk6yDL4ZvfsuJnsG48RmZ1WgE6h9UKWucFBGmdIkSuYMCgmIRW5nZvZetX85T9s1TZGwNj8dzsAk+1aaZaz6VaHUi1OnR3e+lcDvOMBp4DcEow1pLNRjuWotmMEs4Z9+SGYkgpy4BE+ne+SoPWGoPBoHwfUkq3VKvcZy+EQLPZbEsp25zzI1brT/a1+jGu8nek5l8STPzhsT373xNS3n1/9e5HRs/u8Ny+ZJD2TjHO99bJ7FShAqN04eqgt3FqCrvphIYWzYvXTYVHCdNF8SGl+l9QSn3l/OLR1Xfu3rTTJDQ9PpDjV1+/1Pvxj53/utZqHf3sei7wcyyOn4G1M4I53yIjNLiMHFvOGphcwZgCGigIBFFEC3C8UAmwpXWD4BzWUtbisIzDWO6YbAxQ1sAYN3jP8gyCczSSBnjhBeSkiTmYBJixhTqQLRZUtZslgcM49/MCTiwwbpIUKizxrIWDxxgl0eL3KKEUPyirxmKB1VhntMQZoBlJHtliObZQbij+QpAedYSkn2cIUis6L601YDSMyqFVBpXn0Covuh4URAQOwzi2O9tbvZXN38+6+F804mv9XEc9lZ/qquxYB+knFewnNHDWAAsAWnDEw4YUURwnMVrtNqLIsQellCXMRoHTGCcyu729DaUU0jQd3l/SDhbN87wko6RpWj5Go9GgzjeClPuAZJ815oTOs29Ks+yHhM6+GKv4fz2x98Cla+srax+Fe8cak2irzzAumnWBf5TEzjB6UA+/VT3GpAoJVb8XIhd+YvI6oshIeSHL8+/kOX8PwN1pEpoeH9jxK6+9YwC8/yPPPf3rIuvf1mbw8zaOPyniZN6yYrtfabdegx3L6Vxw6EJzDQwlO83ppAoIS1I4xdjFMlhmdthh3LmjFiIHyI1LOIwxGG0caUAwp+3GGCw4wAxZ5xUdlQDjtpTGMYVGm7WsmNHYgrXmzX5MYbMwBn/3kEXnwQQU3Uxgx812ftUyDM3KdiwZ3Hk0RTLaESNVMFo7ZW3jvJOUdou9qbYwXKKbZvntG0vvbGz032aQUQb29BbyZ3LgMwr4pAUOA2gX9w4jMgF9NZtNtJpNSOkgSfpTa41er4fBYFDOptI0RZ7nQ8HJd/30hTGLbXskSVJ2U0PCmZw3uBBHmIwWdZ6dHeTZt9vM/OPje/b/nojkjScdojPGRNaYRSZkfD/zmXFHlU1DFRxX1TFV2HiPfB5/ebUk4kTRwTxLv1vq/PefXjiyfGnplpkmoenxAcNzl5Z/9Lmn/6NKe1ucq7/V0/rb42bjsGTcJSKdg0EA3MJwjty6Np5oyi7oue6Bbp9iEuRgr2IMwx2fuVjh4RDMwrLCHLyI4qlxVbbiHIwDkvFi78fBasroEu4yjHyQnKI0rEtcRCM3ZC9pXGfnEgfH/SL293jF7CBvrnHy8pcFys7Q6cTZ4RmQcmrYuXb7P5k2SLVGrhlyy5FmCsur6507G33dBb5ZQb2YA0ctcBrAHE3AfO26UhOMElCrhSRJygAzGAyQFc6uWZaVSYc8kQCUiYq+T4m50WgMVdLGGERRdM/z+9JOUkrBGDtkhJxPs/SwVelTkTG/enLfwsX315bSJ7gTEsbaWQsrJrlmqLMM4bmw8KnThatSSRiXYOqu2aoZU5iMOOcSUXQuTfPv4Epd/EbqhqZJ6EM8fu2NS5s/8tzTX1PpoMOFvZ2x/hdMkpySknMJ5mjcRdUMUXi3BtI1ZaUIC245hBXg1mm0GSfk7ZQWdCGRw2l2RPs7xRBfO8KCtRaKMZfAeFS4ldqdoF90KLaYHGnrOhdt3NhHMzdTgmWFLA/chu59VKfu/YWGZcM3enkKDGnnFaZ0JYRnYH3atXYdkEtCFqkGDJNQnGFlYwM37q7Hm8BzBoiscwqPQmyfnp86HZr3NBoNSCnL2U6e5xgMBkjTdMhCmpIWfSVJUj6mEAJ5niPP8yFNNN8OwCczhNdDWVkL0eDN1gWt8p+zWX7CZPYfnth78LVr68vbT2QSspZba5OiMhoLk4X3xyTQ2Sjn1Cp1bK9Lm3huVKVlVyYjGR3I0+y7I5X/+2kSmh6PsiPq/shzT/+ZUfmGyPVVZft/zTYa5yxjbaMs4kiAcQalNTjZNRTBqFzALOYsnHMYYV0SgjOys7YgpzFWWBhZMFNAAXxHiXpoz6hUYUgLTyPX2nBwmLLSdBTmks5cwHLUgTgozlJAHB4K7aKaZLw6uIQ4P/OUsq0xjuhhfSac+8pLOM5CWQ4FjkwDm70ebi6tYa2v2qUKQ5AAQyyfMYYoitBqtRBFEQCg0+mUHQ99Pn7SCbsYmhlRIPP/HkVRSVhgjCGO46F/78N4w4nZC8AyOqqt/UGj1D6m8D+e2HfwlWtry0/inMi5gwTIbl2yGdXtVF5nI5SyR/3ObmdHI5MQ55JJ+VSWZ992et/C2++tLa1Nk9D0eFSJSAG4/MPPnPklNhi8q03v522c/DnF+QGbG0QW0LDgxJgqqMYuKBa200LACgGrNbgwBWuOw2388MLHyA4PRu3OIJbxnSTEC8zLFlRqoQELDW55scHkIDdtCyVr5gxed6AxVs50YC2s1sVMabyLZR0t1q9Oq4KtS86mNKArDepU7tQU8twtoxqDLDdItYUCxyDPsbq5jbsrW1jb6EAVjDQ3kzP3JD0fSqMuSCmFLHMW4mTTzsvF3eHkQ12ML7gZUnspORFzjiA8SkI+waGKFhy+ZhHF+63Qn81zNYc8/3+f2HfwS9fWlp+0StsWI01bFfDD3Z5RycP/fb/4qvIJCpPRqMecdCbkP+89iSiK9muVf6dS+e8AmCah6fFoj3/51rtLP/rsU78HlW5Kbn42Y/ZzqeTHDawQwsIYTVeyd8M56R+jtQt4XIBHBtZKGM7BDXdOr0yAc3OP2nBpClbMk9yN5t1kbqRUUKP1jmodQ0Fe8DbAPfiMkb6bdQujPvNo1E0e/mkCiwsf8/cPl3h0IcFTLKVal4SUoj0gjVQbpMZBcTkMNjo9XL+zgo3tFNo6lmFubGGlzsFdNrrHRI/Ya3meDwXAKIrKGU9INPDpuTtFhC07IABlwvHhN0p8NGeiuRD5SPnnwtcoM2bn87aMzWmLT6UqbwsrWqf2L/zO1dWlO09MG8RgAZb7ulZ1ncdu5jejOplx86H73U0Ku1j/sTjnsRHinDLm+TMHDl95d+V2b5qEpsejnRO9eXn7Jz52/stKZUuJ5G+kufqp3IpzBpgVnBW7NY4c4Kp/CWscdVpGEYwQEBCw2kAICcsds00IAW53EpDxEkN4I5hyDOQnh0LrrpxBBUhJQYQo9VKJPMA4GLMVS7bVkMY9SaikzNmSzl0Fw1hroIxx5APfqls5QoIBkOUK/VzBcIlcWyxvbODO8ho6vYHbZxLFzpNx8y4nbbRDf/c7MUoWdN6iKEKSJOUCqp8QwoVKH6LTRfFAiSZNU2it0Wg0yvdASc1PSvT7fgKqWqg0nn0F47xlo+iFgVb/RaKNOr1/4d+9t7q0/ISkIQsgtdbYUQmmKomE3wu7pUl05yZ9znHwW/icPvtxpxuKF3Safk5p/SU4l+dpEpoej/b45dfeyQG8/ePPnd80ae+iEtnfkM34m1mSHDZGQ2mFOBIQgiFXCsYwSCEKd1INYwSsNEUmkUW3UuzTWNzbCRWdDxc+DYHI3halyqqjHIQKQvfeoGTdbcunvgda8yvWkYmJVSWcnYTkC5Nq43Z+tLEu8VgLC45BPiiYcMr5DWmLzW4XKxvr2Or1oU3xPIbBclY2d1wUszRjK2dRBLURMcGf2VQloargFRqy0XNQgiJ4L1RbYFXwqvdc/veG4R+RWLBnBnn285yxztmDi//xyvLdx16zjDFmAHQA6AdhqYU/ryIajOtyqggMD9oV0fVSKJ7MaoaPWauPALjxUY93fBryH9/jV95457ZImr8njfhvRaZ/qdfpXDFMZDxqIFUWvUHuNNMKlprSGmkBEeV5jlxlyPOs+Hvhk6Pv/dLWQVeadmzof6wQUYVPgbbUlHhfwdzEWDBDyWd0EAi//KQy6ovsuHWhSp4rRzowxkIZ999pnqGf5ciMRaYsDCQMk9js9nF7ZRUr630MMrdaS3RBxpzyt+DDFHBaMPXJBlEUodFooNVqoVnsBvkzHz/J1M4Agp/Tv/O7GN+IrYrc4MN+o35ePjbnTUTR8wOj/o7W+s89tXCo+dgnIc4VZ2wT1upxzLf7PUZ15Q+S8EYty4Ykk7JbYuyQMursUwcPt6ad0PT4UI9ff+Pi9o8+d/7PjM7XpMneVL3BT6dCPCdiudiImsiths4VpHDwkeCshMSMcSoHQkgIYcC5rp1XMMbALQ9mN1TphZBPWLuM2ki3YxPRqBvWwFS6VlJ3AjgVCKVVuROUawWdaaRaoZ9pMMGhYNHPFLZ6A9xdW8PKehe9vDDbE06x20kG8doESdUqQW6tVqskJ4Q03nDmVgfb1HniECnBJx/4X6Oq75AtR89DSgxOnYLPGCE+0VfZ32gBa08vHn790t3bj+2CJGNMM8Y3LKBYTRGzG4HS8DyNY8ftZp/ofjuioQVWIeZNrj6utf7djzokN01CT8Dxa2+8owC8+8PPnltnSr/ZlPK7MmW+p5+nz3CBfZxZSMMguZvLCOaq+0gwcHBom0NYNwPS1pTVsixZVnooKQ1V6dhhu+0cOkTfhpLR8M06GTs73M3YESI1lYw4RR2TBnJroAprcGUUVK6htUVmAGUZ0oHG2tYWNre3sdVLsd7tIVUAl4WCBBMYnn+5fSNthoMEJZwkSRDHcbmUGgYjf49n1OwgZEn531NK3ROcqIAYNyQP4Tl/Bjh0nrnYn3P9uV4+uN4C/gEeglnfB5iFFGN8wxqtLB8N5+6m86mD5HYLy1V9xlUQdNXvVWndMS7aBup5Y/ReAEvTJDQ9HovjX755cf2Hn7vwlWxgLqs8+13N1E/w2eb3cClPWM5aGoW1ggvdMNpCcA4mBIQxEEUwKgNSsAw5BNkwT/CNjbFNLkdGVcGgfrei6u91nZAP1zkL8kLOSBdeRIUtt8qNU8c2BgoSAwUsr2/izvIytvsDKMsw0E6FghfMMUNaRmDOMqJQ3YZnJ05JgGY/xFALu486/bG68+cnIUo8QojSFZeSnw+z+f+2rkr3JWGqkl2ZkER0JNPpj0idXz17YOFfXllZejwDHmMKFhuwNq8iudxPMqqya5h0J6iu+5mEeFPXBQXdUGQ5O26sOQrgnWkSmh6PTyJ6420LYPmHzj+1zjS7aTf7fziQ5qdEq/HNUsaHJWfCAGDKwnINzS2EtTCMQXMOYS2EMZBCwHAGzvgQhGQLmjLnAihcVst7zEk27NyERdIxdCPae6tMp87AK3Fxv+uhGUj4e7rQjqOfaU+KRxkDY1BAcBa6sGPIlUKeKwxUipVOH8vrG9jY6iMHA2IBQMBaQEEUGnjaGfBxViguWDi7Jl44xg4rI9CO0DhjtXFUYV+FwZ8BJUlSasyFs6KRxUBFUPPPZfhaS2adlKcGWv91qfX7Ty8c/tKlpdvdx+26v7O1ls/JZNNapFXdzKTdyyTd+G66ofD87nauVPXYVGxoxvbnWp89ffDwH7+3fLszTULT47E6fuOdywrA+z/09JkV5PkltpV9S58Pvkc2kxdk0jgiBG/CWgirnfp2kQiKTT/Xn1jm7COUhWC8pPy6qrtIRsw4DbsQNuA7q+shJn8Pjdp7XvrT5TRbWc1aOJlsyyxyrRxzrVAQ9+c+xhgYcGTKIFXO2E5rg36eI0tzbKcZbi1voNNPkVnACmdVoS0D44UShVLO94gLSM7c0i1IbsglIepEKBFRAvITQ7jIWCdqGeyElOw3/7zFcYxerzdUHPhQ6biKe1Syqk6WPIZkz/RV/rcYY3fPHTr6ZxfvPI52AqwDa7ujoLVHlXzq/s1D7v7mMp0/H2vVhmMGTpPQ9HgMk9Gld7sA/uwLT595hyv12/mWupDKre9u7Gn/oOT2Kc4sjBCwrNAVMwaGcycDVAQ1KQUk4xAG4EKDa/enFKIwvUMplOo6IIAVi0q+kHUVLBHOeMh2oQC/diA2WsQtzOiscbblmgKMUrBGwWoDbciMzkJphsxY5EwiB0M3zbHVTbGyto7VjQ4UZ9CWwUrp3oRlhWaehtEWkruEpHMFZQoBUcahjYGUOxAlwXC+IZ3PlKvzsJkkkPkdUZ7nJSHBd1j1YdJJJGX8f+8nO4L3qMvy5J/mcqhv6WWDn+RcrAK49vghcqJjjd0EoBhjskqoNLz2qhaD6+ZAu+2gRi3LjuqYqu4P/9oRJUxsmobnZ402s/gIa8lNk9BH5PjNS+/24QbLV7/3xIl3BndW35vZP/NfIRKntNYw3lzD37FxAQvQ3EJqBi5ckOaCwQinP8fhoDfXHPDC6gHln85TbljUyxYPvGPJzbzOx++EKOG4hVKigbvZD4M2xRxLp2BawWgFFLI8qtB/G1iOvtLY6PdxZ2UNG9s9KGOhCy8l678wD1p0QmTOdZZ5AURICV5AhNQBERkhFBWtCz6TBjQfGvMN7nwYLuyC6iC/UYSFKvLDPYSFODmksvSHcp2/em7xyL+5ePfWxuOVhFifA6vWmgzgcqh7nlAr7vFLrPdeM977kJaxI9bqgwAuT5PQ9Hhijn977dp737144D92l1e/Wy7uP2aZLW5Yx46zHimBspDlHIbn4Fo4GE5z6CAACsYBblxS4swZ7xWjoXv+9MzmHCTnqN6OPu4UrlHAa6YQHVVF0trZ8mcwljlJHp2D6RzWaFiri3/HoJnEZqeP26ubWN3uI7UWmXZq3s6Zb/S5CjfWafmUc16ayjUaDSRJUjmXeVgBzw9AWu+wFf35U9V2f11XFCai8LWGBIUyiEfxyUyrn4uUvnbh0LE/fvvOjezxCdg8A9iSNSZngt8L49ZAovfb6UwCzU0K5VURG0Yx5sr3wPm8sebwUwuH48tLt7OPYryaJqGP6GEstiMhMs5hOJdO7sdYKJOBWQ5GHQ6nQEVzB11CUFQll4PSQGxz3A1HyceJm967hIrCxM/BcWRGFzLhiufQClZrsKG9IQcGRpGEhcZ2Zl03xQBTdGZsTPVJhy8w2mg0hoRH/T2gOhLC/SaeENIjKwdf2idUVRjXcY1Sah4XkLkQDW3NC301+GnmIKBLj8s1zTnLOGO3tTEZ47bWI6jqv6sSwSg4c9Q5rYKeH+R6qFJN2ElCYlbn2dNG6yaAaRKaHk/O0e0PDszPJEdFJGMBOPdTkjAoKMi2sODWcOQDy3kJ25kiEYFYc2xYAaCuih++aS1co7Gjk+V4CrpMSgACpQQnRLojxVNQlY1LQBxeMGUukclEQsQxgLSQDALAnXI4G1Np+ppsftCnOVC4O+UH9oc1iPYTDqlyhwlkEghuXIKpkvqp1J7j4kBmzPdxlV5++uDhX7q0fPv2Y9IJ5QzsDqxNRyWIcWsAk0Cau+2A6iDRUc9bBcve83yMtYy155TWbQCbH8VYNU1CH8HjXDxz4tp251sa++OTbgavwZiGZLxgtbHC/8eAWQ6jNMAdvMUg7pGU4VKWSSiUmhnl5+L+HDaiC5MQJR7HfNNg1kCjcMiDLVQb3LSIl2KiReAAg2Ucaa+Lfr8HBiCOgdQKGBRzjgI2rAsmxAYkBhztABEMFnYp4wLaqGp5HCxIXVee5/dI7tzPc4VqzeGAvqqrKof5XBwfKPVXeZ5eP7d49N9dvHtz40NPQpzljPEVa1VWf73Vewvd71Lq/cB0u+mARu2OgbGGBk5rrfcCuDVNQtPjsT5OzRyQ3U739K2s84Mx8J8h4vthDQANZp0xnWQM4AWpoDAiBQBtTWETZEsHV6MBCwFhLYC8Ft4ZRY811n05g1VbaNCZUgrIT0KOwGCdE6thADOIpHudEAwCw89rmIWARRLFmGu1sbyxBZUBGTQgi0XTMQHbp16TCravAUcuqZMw0sYFnDoTNJoD+YGySlbJf5zdVOn+4moIBYaOsd7rFAZ4updl/znnYuX84WNffef2jQ9VPoYx5JyxjjUmCxPPB6knt1uq9qjCo66Druq0iy8Ozhcs7GEAb0yT0PR4bI/Drf0zdzvrn+xD/20GfFYA+/NcCQpCzGgAzg3VAWQFM0wWA2rjgpH2PIWsZQAMdF5YKhgnaEp/Otac06yrJCgUSagMcEMdkWeJzO0OzFZ49zDBAAgIGDDm2HXlQmx5E1swGLTjGHPtJiK2BWXh5IiiBCon2ne1JBrnvGS9EQOOnE1tYW5njCk7E4yA9qq+txsVZ98ML2TF+RX8pDDgJPtBlJz8n9N755xDc97SwMcHOvvPRS465w8f/7N3bl/PP6xrfGl7zcyJRtdaZKEdwigNuQeFT8cRCD74DpDPK2XOHN+70Ly+vtSfJqHp8dgdC419h9d6Gz+YQv9dAKcioL1nTmB2pgUOC2YdzAXXUJQBHOCFZE2RlBgJIpChHYdhLohz5mSliXRtYAuJGzgx0TqWHGOeuZCjQnNaPAJ5GnHn5sr8ZOEen1vjkggrbCV2QigK/wVIyTDXbmL/HoHlroZSFlZpCM7dv/XsKyjQUudDAZ/mP9ba0svHWoskScrZiVKqlNRJkmSIVFAHDY2i4FIAlVIiTdNSLSHP8yFYsKrK95PGPbpjNcyrKoWG0CzQ78wKKHZew77UywdrLeB/APDmh9sNsS6AjrXWMMZ4nb8U4Par/Pe0owgyLPA6ivhRB3c+CNNukmJiaKGZsZlMZU9LkcwAmCah6fH4HCfnj0a9XvepjcHGz2YwPwzglBCIuAaEKIzQYIdiNyUIP5SbMilRt8JgmYPFyhrcmsIjyGFrws9VpcYcKv50CWc4GBvHa2POocglSF+rzoBb98pY2cWYMjGWUBoKnM9oCGsRyRhW91EqCDHm8pc308myDEmSoNFoQCmFmZkZxHEMrXUZ+ImdRsGKkkSapmXy8nd57rdipkBECU5rXdKxJ50FjXvscfI+dSKcQ91XFC/kZvB93bS3evbAoX9wZeXO1Q/rmueM9zmwCViNEVY0D3LuJoHdHnQeNEkH64mZNpW1p4zWH0lbh2kSekKPE3uOzna7nee38+3/NIf5ThnJYzRX0ABiKSE5nNIADfeLAF7CYkXn4d+uhrlAz2CGAj6lkyp1BIy8GdmY79oi0XAv0Rj3GpkJNFH5zmtiBhZOC09rBQGgFceA6YMz0rMDuOBuwbUIHO12u+yAoigCAKRpWkJvnHO0221kWVYqFxBJQSk11AWNEysdB+0QHEYLqpSIfHr4/SSZcYZroe2EL3Tqw3H+6xVxcixPBz/RTfsbZw8e+adXlm/d/FA6Ic5SDqxbaxWAyD+voeVGaMsxaXKeNBHd7+/UfZ5VO2jFV2wZDllr9nwUY9nU1O5JTED7Tsz3Br1v6ar+/x5CfG+j2TgmZQzGBQRjkABiGUFKknvZxQXhw2LMFN3QzpdgFoLZe/4++ssGX0UHVNHpuO+F0Jy7VO09iawwe4OBFBytZqPQxKNcZqFyVe7+0MyHKNAkh7Nnzx7s3bsXURQhyzL0+/0yGRCEE8cxmk3n/TYYDHatll11+PMYfzbkJ6FRlPhRVOw6CaGQdReyHavsPIiyLuLkZM7sXxtk/e99evHogQ8lYHGeM8bWYaFGeVH55/SDIi3UdcAP8ny1e12czzOGfacPHP7IxexpJ/SEHacOnJzvD/rfmiH/edlKvpULvs9YRzgQXIBbJ7jGOdsZ9lvc09VUdURDiWiim2+CmwpsGP8LHyP4kfXqIuYRCiwAy3jQjwGcOaVuKTmiiINz9z3AgguBSHDYIlkRCy6KIjSbTTSbTTQaDRw9ehT79u3D3bt3cefOnaHOhMzg6N9prcskFNorhNv645Yl/Y4jjuOyEwltwh8EihtXmYeKCf6icJjMhBACSXwmzbK/zQb9zrlDx7548c6N1UfcCeWMsXVjjOIBZT7s5Op2dh4WVPewmXMjkxLnM5bZRWttAx8xk7tpEnqCjrOLZ5qDQf9jiuv/rDHX/rQQYh6wzksn15ARh1UMzKRuHGIMCpU31DHEHufDgpcdkeu3qHUvnFC9XSOnJ6dLV1lrHauOcwHGOGZmZkoCgjEG586dw+c+9znMzc2h3W6DMYZms4nBYIAvfelLeOWVV7CxsVEGrDzPIYQoiQM0N/KN5uoMzsZZPzPGSoiPpIKIIj6ODj5Ksid8jlEuoD71O3wPw9+XiYnZM7nK/4ssz/T5w8f/wzu3rz+yRMQYV5zxdcDkk3Qf/jLubpxXH5aY6W6SzyhJKC5ECxbHYM00CU2PD+/QKj+qbP4zUaPx6TiJ5zl37UjMAKU0wCx0FjkVASnBOAfj2LFwqICzipAe3roVMNjuacKTdD7lM5bCop5RXMnFw44cj4cjk9q2ZRbacORZVi7HMlEohEcRZtrNcq7DOcfzzz+PZ599Fmtra+j1eojjGO12GwsLC9i7dy+ef/55xHGMV199FXfv3i2lVKiKbjQa6HQ6I9WzJwk+4WyGmGrj5kGTVM+TBMyqRERBu87mvPi9lmHshYHK/0szMObcoWO/d/HOjbVHlIUU43zDKJWHs6txAX6Sa3ZcB7nbBPWwCAyM84bR+pi1Np7CcdPjQzmeWjg50+t1vklL9tlmEu8XkQBnDAwWlllY7tQPuI2gI4k0V+jngIwYJBikdR5AsLYI3hpgomTDBdmJADBYpmFNwVQrA64dmjN9UHC7YR40yFwfZH2DPcAJqjLhxFCtca9dMEgZIZIJGo2kTD5JkuDgwYOYn5/H1tZWGfCTJMGBAwcwPz8PzjkOHDiALMtw+/ZtrKysDAmKEqzn05jDrmU3UEuoHRfOMybtqMYlojC4jkpEPlTnz63oT601wFjbCPnxQZ79lyxj+flDx770zp0bGx98DmKaM74Ji3xcsr9fZe2HTVyYlKU45o0n2phDxphkmoSmx4dy5Ong0CDrf0E22kdZsW9jAYhIwjAgFhxGZ0iiBAotbPY62EiBKG6iZQcwJkckChVtBmhYCOZgLg7uugcSFYUAYwbGU0nYuaHDLEBZq1ou1Fa3WvccO3MoM/SPOSsWZcELejkFlaKXM9hxexUCxjo1CBknENGOHTfgqNbz8/PYs2cPOp0O+v1+KZWTJEkJu83OzmJxcRH79u0ryQq+n4+fiIjdFu6a1CWEKoO7kNE1ShduN0lolPX0pEkzhO/8pGuMaWvYF/t59l8jgzl36NgfXbxzY/2DvhWssV1WiHn63RCprxNzkSj5vjpEnf7fbs7x/cJ1k8KofvKna0JrHVngoLVof9Ri25Qd9yR0QQeOJVk2eNFK9s1RFLU5BQPOYUn7gO2wvRqNFlrtOWx2+9ju5bAiAoSEMha51lDFPgq0LeR7XHJxCgk7dtwWjuocbu67hMTKr4myzP31QuUNyq3ZYcwZC2N02ckYOEdVwEJyOJO+KEKr1UIcxUOkAhq4SylLujaZvFGyMcYgy7IygFH178v30EIrfT80V9vNfIBmQcSMo87tA+okhl5j1Vfo5lr1VcodxckMT5JP9E32C2mWvnT+8LH9H+S9cHdrVcGiZwFVlzz8hBkG+kk+l8fFjyiAejk43wOG+WknND0e+aGUms+s+u6o2Tgk5bCQKIoEBCYguIPZZJxAiAidrQ10swzdTGJv0gCgEXHpgnmhKGCNk8wxVrtxDFkgMAZufaVl7nVCbOR2/kO8DZ2unAPF3XcsvUb3/FpbcCFLeFDGQNxswEYSkZSI4mFXUq01Go0G9u7dC601ZmZmIKVEnufodrvY2NiAtRb9fh/dbrdkyNF7JHkdonpTQC4VBnbBavMfM8syKKWG7MMf5LxWESQmITqMgw79Kr0sEISctbH9RC9N/w8sY//D+cPHfu+d2zc+OCdQy/rwbA0msXCY9H1PMt/7sJKRAWaNtfOnDh6Jry7f+sjYOkyT0BORhLITCvqbGkky6wKuPxAvwnFBX2akIiAFRJwgMwZ9bbEnaiGJGJhWiJhF1u+iGcfIstTpyTHAWAYLU7AHiqRjLSx4qVwddj2j46R9wC7JvQ5YOBM+7GB7lIRM4YVkYZFnyu1JRTFM5IgIggv4sE2328X29jYWFxcRxzGOHDmCZrOJW7duYX19HWtraxgMBlheXsbq6mrJgqODuiH/76R0ME5YtC5ZUOdlrUWz2bzvZcdRVgUPo/IPjfAoKblIEs0A7IVenv0CFJoXjhz/nbdvXb/1wQRlpACyqrmXryO3Y45odwWlfVgJaJxXFeOspY05aq1N8BHyFpomocf8OHPwSLvb7zzDY7nIpFMFZQyekoCDxlihii24hLUG2mok7TaytIeuMljv5zg+ewDC5IiZRkNKSGuQSIFcKShroY117qZUORaW3MbT4WGsqrqsS0C++dx9Fr1B8DClLwTp0QloY6HBkCoDISUABs4ZoihG6exawF4bGxu4fPky2u02Lly4gEajUXYvWZZhMBhgaWkJN2/exPr6+lDg9TXWKPlUVdu77WCstVBKDfka3e8cKOwOwi7ofkkOVQQG6iy9TrOlOXsu1eq/ttmgfe7Q0X998c7Naw+/P2Y5gNzXjwup5H5CqusQP+xj3Czu3oTEWkqrI8bYBMD2NAlNj0fTBel8n+b223kj2gPuMlB5gRbQFCzASLa6UCE12kBGEiaX2Oyl6A8G2Du/H4fm5xHrDFHSRNbfRqPRxCBNoaxGriyUsTtzDlVUk1rvaNCxHZ04BlaRX0LCwoNWh064lIHBGjsk40NJyTAOWcy8ZBxD7fRJOyrfO9Ambt++jSRJMDs7i62tLcRxjG63i8FggK2tLVy7dg1LS0tDMyI/MHDOS9WFOhho0oo7DJRSyon//W4TUl2lX0dYqNspCt+jP4ORMkoU2Pl+lv4dnZmZpxeP/moUR+++ef3qw4v+DDncTGhndQyj3VQfJ3htN0lq6P1wlhjYRWNM9FGKcdMk9Dh3QQtHeb/fOasl/lwUxzMoCQnM2R/QfcW5SzzWOO8exgDugjKPG9AW6A36eO/GLRxe+DhaookEGraRgLEcMoqgrIE2cElIaWSZgs40tDXItYLRCsY4nbbCeKika9t7ULcHheGGIw6NIBjCIbpj9cXNNqzm6HZSZCKCTDikjGCsAedRsbjKhgL/tWvX0O/3Sw8hSjSDwQDr6+ulqjXBbARBhfYBo7TbJjlCBWvqKj7IanuSLf5JF2VDP6KCLBLZKD6Xqfw/NWnvQNs2/8mzx05efPPG++lDgq0UAxSsNTZIln5S91lz/n8/SGJ/mG66o5Jk9fOw2MLus9Z8pHaFpknosa6EzD7NzHeKOD62A3mgHMyzgBbN4GwVyD0VtvClaQlkFljd6uLNi1fwqecvoDUzA6Hb0KqHJhS0MdDWQhsgS3NYy2AU0B/0oY2G1qoQ8MwLoU3lGdJZGOtX9MPSOkP2EGOD3/DvOviNZlIcnDkjOiEluIwAESNpz4JlFls9A9FUSIQEYwKc8RKm9AM9Ywy9Xg9vvfUW8jwvf5YkCZpNt9hK0jlETAgr/jqPodCEblwCCmRxJmZw7SZg7mYoX9U1VdkP1NmOe++fa85Pqyz9qa4aHGwz/KNnjp547a2b1zYe+L1xpq3z3r1n97lKA2/Sc/CgWoAPvfMJPgNrrbTAHriZ0DQJTY8P9ji7eCzJsv7zEOK7oijZyxkJWrKiz7CFvYIouhJbQk9gDsDijlEDbQxYHCOREm9dehfHFhdxcP9ZNCWD0QkYXFLhQkBrg3SQQWvAaoZmqw1tnBKB01PLkecZVJ5DaQ1r3HBe6RxKaUedto5CrZQqhsPDy6334t3DytL+zwQX4OUXgxRurydOGhBJDBY1wWQCpAYGQDNpDPvs2HsZT8RkazQaQxbepKpA3/MTF9GxKSAQVOcnjlH20XV/+irWPjX7QeG4OgvvqoDsKyXQZxBCbX43UdcFVqlH8EbzqM6zH9jO+0dbNv4H548c/6qQ4sab1+4fnuOMaQsYa62tUp8ulb+FGHr9ROmvSy6TKF5MokYxrnscLYuEez4bb3eIW9hZxtCcJqHp8QEnoONMq/xpzexf5VH8NOc8Ypw52K3Y4ym7BeYHeDYU0gkUE0K4xACNPQuLuHT9Bg4c3I/TRw5iZmY/hM2QZyniyFGVZ2cEslQjSxW44OinHdcZFYFYqRzG7OzNGGugFSUhA20U8jxDluVlxzQ8V+Fe0HZwHnU6gnNwwctZkBQxJBcQkkFwUXQpEeKkCREnMDyCljF6a1sQApBxAguGOI5gjAYT4l71bS9w+UZnoQ6cb39NxAGy/KZOqGqHyv+3owKPT3bwFbsngWoedmVeZQFe9XP/nPnVexVNukxmcbLfSvltvSxbiHP9L5to/Otnjp+8/Nb19zfvs8uzDFBV3MwQkqvr7p7Eo7h3Wox9tBZWp0noMTvOLBxjKs+eykz2V20kvlvGyX7GGRhncHmIO900a2EZA4MphD5RyhMwO0wa4FyCSwaTGWjGsbzdwft3l5A0Ypw9cQRJHANcuEVP4eDmJGFQuUGW5+ARczbdlIRocVNrGBgYq6FyVQZqW3RCeZ4XgW0InNtJk2QjDrc0OwyjUKISEJwj4hxC8B0l7LgBESXQIoKVDSxt9SEEoI1FJJwAKCnmVTHCws4lhG+qfHWo66EOL4qiSgvuUVTpMDhSsvJFS4eoz8B9s9p2C9vVEREeVMHB2bXLto3Zx7I8O5APut+U8OifPH3o6B/LOLr+1rWru1LX5YwZBuQA7KgOkBZq69xtH8aM6EE61Ek+j3s6IsEbYNj71OIRdvnuLftRiHnTJPQYHacPHGln6eBMqtOfMpL/RCNuHebOmwCM5HWKQM7YsCippf9n916XWuUQjIGLCJYDFjEuXb+JXjpA3Ehw+ugi2rNz0P0eZtrNYmfFQEYCUkfQpgFbwBm+zUE5VIdBlmZD3wND2QUNBzS3UGsoADNedHPF3AdOdJUxUc5JOGeImYCQHFIIRHEEGTcgRAwbN7DRz5ErAy4cbGeZm+VESVwbBPxqnv67Cpv3bQ1IWSHP83JJtUphIEwikwQzX7JnEp2xUXBbVaB8lNRkX4zV75QYY4xH8RHN8j1dlZ2NM/Vvmha/cuHYiTffvnFte/LHZ4YDg1GyRPQ6iG04rpN8GPOgh724XT0jYom1Zo+1NsJHZFdomoQeg+PU/mMzSmWHer3ONylmftRK8ZkoaSwKITinwMy4+9PrKFgIv3HXZXC7s0tkAXCrwbhwigg8Rq4NVrt99N6/gUGvD/npb8EL508jyxUA5rTWOIPSQFO2oAs6sr/8p7V2ZISC0k2uo/5NQ/Mh6njo9wmCs3AeSATFESlh579pTsIQF91RJBh4JCBlDCsi2LiJjtqGAYPlHFy4GdkkSYCSnJ8IRlXNNAvKsmxIviacY4Vw1aSBexTUNsqraFI6eN2/qbP5HjfHCOHNUWKo/nlhUdy2Mnomz9L9Kut+vKHj/9+5w8e+IqS8+db18V0Rc51Q3zeuH77uTMlsrIIOw2vjfhLQbpLYqG5o1ztlsIk2Zs6aaRKaHg94nDtypqGUms3S9NB2d+Njuck/rxk+HTebx+MkmYmiqJyfcFbAcUU/5DoGu0Mi4ztA1zBXDiAdBRiD3BhImTiSQiOCGfTx3q1b+P0v/QFmY4FThxZgjQIXgGUMYAZCcgge11Zo1u4MtktigjHQ2hTLnGZIWDKkzxJcUgU9FHsnACwkGUowCyY4OCS0lMgsgxASm1ubOwu7UiCJYyhrRmDrbGQwCtWkqQMaDAalyV3ofno/VgK+YKU/O6t6DQ/a0YyiXY+C5argwCqrh/B7VY/pw50iihesMH8+NeqIVen/klj7r545euLtt25eWx/zPjQHUjsiyPvXGl17DwtSe5idTt33RnzOsTF6j7EfnV2haRJ6xMeFY2cTWLtooV+0PP/Wnu5+U0+n5+NGY38SRTOkHeZX2ow5M+wyUBcq2juLQnZ4M4f57qQW1upiqO/UEZgQUFZByBgyaeLqrdv4D1/6Mv7CS5/Ggfm2s8k2gBAc1mrAFvMZRnINxRJpsSDLuQCshTYGMMZBd57hnDa6DAZD4pIMDo7D8M4Rg7OdYEwUo2cLUbABGYyzpACH5e7na+sbePXVr0PICMzTchPCyfmwXQYGn0XnEwgGgwHSNC3nDX4SmjT5hNTpKiZamOgncUh90LlGVaKp6pCqXl9dh+kngfDflwmL86a14tk0zw4O0u63NYT85acXj/yOjOT7b924VrlXVIwYB0ClTVYlUSI8/w/iFfRBJ666RFRoN0ba6vmP0sLqNAk9ygR09Mw+rbJnIe1fymE/ZyN5HHG8N+Zc0l5K1RcF7J0VmkIBwAZiixTACR6Bg8CYACwvgr82gOXghgFMALIBJBZvvn8Te/a+jQtPncSFMycQMQZuDGIZQcM4jTbLAM7AGYc1xfM40TmXKBhzZnJ8x9rBlpp05UssCQOWofi38LgKRRVd9HHKAEIyGKPArYHgLgQpaKDojzY7Xbx37Rbae/eDe2Z+DLYyCfgLon5gIgjHp2RTohkMBqW+G/1OyKa732A2ym5hVOW8G1WESSvvSY3f6joq3xbctyaoSlp+V8SEPGgZmx9ofUKpwacbiP+n84eP/vE7t29u3JuEGBhY6l6KvWeJ2Gc8hrM/3/q7yqZiUvitLoHdL1mhas5X1a0aBglg3riZ0DQJTY/JjvOHT0daq2Nap985sPlPcxY/b5k4AID5N0Vl8vFvPI/aO7z86aZDlrjOflBhLnFol5IQcee5A84BAxgOiKQFDYY/fvNt2Ehiz555HDu4F7GMkA5SCOEqW6dLZ2G1dYnERfqdYErECLbzmnYUtyng7ji9MuaSY5FRdxi3jIFZ69xUwR37zyo332KskBBy1HTBI6Q6B48jKGMhRCHzwwDOWU2tXG1vHcJJ1O3keY40TUuLb9+ltU4x4X4Dke97M2p2UEf/HgX9hYm36t+ME0KddKhfBytWJTCvG4wsFyeVVnu30v5T0uAfPrVw6DcuL91ZCgYjmgE9WJhwrhUQISq/Hwb5h0EmeNjdUdVnUdxH0gJ77LQTmh6THk8tnpgbDLrPGWH+Mo/i7wKLT2iLpi0gKoItQvit6mscnFB9I9iddGB5ucRqwRzFmzNoAKLRQNrv4uXXXkd3axM/8v1/EawhIJIESudIUNicGltAXKTeYL219WEtuVI/wZqdpFkmHAz9t0sttvg7GewBknOXcGDdPKiA7zg4NGO4s7yCldV1J+EjGOI4AeOsZN6xCbsBCvy+ZxCx4TqdTtkF0Swo/JweNOBUfYXBddT7GLUXs9uZ0SSPURfAq6jl4yjfvio3XHM8x+PkRaXyv7fV7y6c2X/wFznn719evmu8smsAzwGxCi4MZ5HjVMbv93N8xHMlYa2dtcBHRrpnmoQ+wOPswWOLWdb79pzpv81k8jERxQegNfIsK6EeYmf5M4Zw4P1gN4tn92C5EwIlGK3oZCzjYCyGMAqDQQ9vvncV27/8q/jrP/PTaMURYsGQ5xlYborXSRCH6zhM+TxFP8Roh8lZF7mU5zum2tJB3BR/J71uMApe9J6dNBAACLBixmRhmYBlEXJtYMChtEUzboAVLA0hRTlfGjUbCKnYpIxNwqX9fh/9fh8AEMfOIG+SxLPbZBDSmcNA7sNcPuy1GzhukmunboZVl0zC36+C3iaR+/HfZwF3RoyxpzOt//ZGv3toNmn9o7P7Fq4YY7q50pGFyQFhxnWVPuFjVCJ61B3QbmDP4HeFBVqYJqHpMep4+tDJhsqz05nu/6CW7K/EzdmzFjtSG7RxL4RAkiRl4vETUZVs/rhEVP09XgqMMgivI6K8wSG4RJaniOImokhi0NnGOzdv4h/9i1/BT/7wF7DQjiGFKDyHjCMIMMfWs5aAuEIuiLqsgjUn2L0KX/4txYukA+t2odw8qKCaAzBWF9CbU9A22sIyDsgIhgnIOIGxgCgIHcYYcCsgizkaoUJVG/6+ioM/J6JqfjAYoNvtlh1QkiRDVO4qFtn9JCDfGsKXBhrXnVR1xKPmUZPOrSahatctANdBXVV096pA69lZuwAVJ0eNED/VU9libNg/klx+3WibWKAxSYJ40C7lw2LPjWBScstYExO8/2kS+sZMPsxodSBLe58wwvwUaySfj6P4KGOM+xbQflU2DoZ7GLABY7yyP4IFLHOzF1YM9LNcgbXa4HmMS9dv4Td/+3fxfS99Mw7tn8dss4VsMIBWOeI4AhiDVTkYEyXw5xhzHM4UDzClzJCfhIrgT9AcTJGnuHMvsm7eZK0BrHLSQ3B7UMYwQEawQiI1BpevXMXrb76FKI5hrUUcx5BxVAZz38G+7sb2uyI6t0op9Pt95Hk+pClH+mMhI243C6R1gdKHj6hDDruQSTXMQkrybiwaJkk+uw3iVXtJdefL7/qKwmy/Yvn39vr9OZYOftPk5pYBjlprRd1r2q2PUNX+1YdhfjdZt8YadpqEpsc90Nvi8bl00Durof6CEexHk9bMuShJ5n11AVrmpABJQ+4QqqjbmblfmKWQc3TYGLwZDQPANCwYkkYD3U4HgksIKaGtACDw5sUr2D/bxMfPP40zJ09A8AgQttgjoqVSB6mZAvgzXvOzM+XxXg/jpegqqYHvCHAzABqwAuBuNsStATiHtQwQDFZK5BbY6vRx7fZtvHf9OuLWPMAFwBmE4MiyvDi391bb4T6OL9FjrR0iIniB8B62VxigQ5rzw2JK3Q/kN4qW/DCo31XBetT36p5rFHOOIFFjDLgQs6aRfLth2UI/776jgSMWaIw6T+MUFUb97qNOQHWzysrvM8TmI6SkPU1CD3g8deikMCo/lGf9l1Lkf81K+fG40VzkUvLwAqJuSCk1xK4ie+gqReCHASWEOzjFqykVfqxRyNKdxVFwDsMMGJdA1MDX/vR1RFJiZn4fFvfPQzAGpXNY65KpLFKQgBMzdcINjp5d/olKRaHy5+61OdzQwEF/HBSIrIPqABgmACbRVwa9TGOQa2TKQnKg1WojyzJEEdGs7UTBWWs9JDWTpin6/f7Q1r2UEkoppyaBYSpw1ePv5rOr2r0ZF+SrElHd7GZc4L0fxYVxjzmKtTfOQ8cnKvjfi6K4mYN93Az6x2HBGOcfSjfwsNTNJ+987jkiY8xHRkl7moQepPtZODaXDXrPaKZ/KGf2h0XSPBnFcZMYVD7Wn+d5KW8jhAAtpfrCmP6sIZwLEU5OrK00TctZRYmf00ykgPjyPHfuqqxY9PRtftgOnUBwBgtdLo7CGEghYJkENwz9LMd//PIruHV3FT/2l76AhflZKG3ABIewxpnGwSWmOEqgjYUxmVseZYAmKR5rHRGBFYHKWrDifVljIYWD4CwshJTI0twRDBhHqjSSZguZNsiUwWanj//5F38J15bXEDcaTmbIaCRJ4lQTivNPiSjUMvODgBACcRxDKYVOp4Nut4s8z0urB9/GmooJP3mFAbRuoTOkDodQEC3F+rYRoyCiSVhzYbIJi5O6/aC67macKsQoqLPq9Y+aP/lW55SUhBC80WofGAwGlarfPtWeYE3fKNCnwdfNtx5Ekud+Elo4H6s7/97PImvszJG9C+LW+pKeJqFvwOPMwvGGUfmRQdr9tGLmp1kUfyKOk0VfCZmGzHnuTOAGg8GQz4k/B/D/XV31RN2S1hppmpbJZzAYlLBelmVDNgSUlCzjsNzRapzIQSHJ73nQ3RsHnDqC5RIsTqAVw6X3buCf//q/wk//2I9i70wDKk8hhQSMghQOmlO5QhTHENLt1xi2M5NinCPigNXOY8haAzDtnGKL2ZAzkstgNYOQEoM8BxcSzdlZ9AYpbNzCdqeHX/zVX8et1TX0BhmsjMBFVLnrA9w77/HnDsR2y7IM29vb2N7eBmMMMzMzlQKlfvDw2XThjK9OFqiKlReSJap+HsKAk3RVo+C4ujnPKHLF/ahnT2oNPi5h+r+3G3HY0GbjSThGQazFjl1krGlZY4XDrqdJ6BvqOH3w6EKe9V/Mob6gOb5TJo3jUZy04zi+Z8CslCoFL6lT8WnY/uLjOEICWQjQhZimKZRSQ7pmFFABlIlKSAHNxivlF6/cBQBTzGmKhVQWt5BbQAiGS1eu4Rf/xa/hJ37oCzi4bwZ9NUCTc6S5g/e4kMgzBQvrYDGBMlhbpWCLvR/OAC4F8iyDlBF44VbqAr9TRLDgsHEE3pjF2nYXygLvXn0Xv/+Vr2B1q4POQMFwp9IgRRQM83k5karF1j1/oO3tbXQ6HTDGkCTJ0GflL49S0qmCl/wq29/aD11ZqZuqCtgE2YbXgz9L9K+JB5kb7RY2ehiQVd2MqM691U8mdG9NOlPzz/+TlIQmOLfSWtMmYsY0CX3DJJ9jidHqRK4G35dz859AyPNRFO8Pg5Vf0ZKytDGmpGL7lXgVDDeK5kr/Lo5j7NmzBzMzM5BSotlsQmuNtbU13L59u4SJHLxj3YC/Zi5jWN0MyfHKTFFqRa0ZmDyFzWPcWFrBK6+/jk++8Cz2zrSRwkBwiZg5SR7GnJK3cSZEjtZNHaCHCBpjEMUxjAVypSDjBFxIZP0+tLXgkUAvB9ZvL+Hu8irWOx3cvLuCO2tbMCJGzgADjphzCMkrGWtVM5eQBZdlGQaDQem2GkVR+flRYgvhG+p2/blFGAj9Ljes5usqdh9i2q0S9266krqgf7/eQXXq43V7RpN0PFUQ4ajk5heB4XsMl1Y/KC2++032u/uMmdDGtKy1fJqEvnG6nzmVp8/nyH/CCP79TEbHGeMJDaypk/GTT7/fLyX/KbD5cEtY5Y7avqeAR3Th+fl5HDp0CIcPH8a+ffvQaDTQ7XZx69YtCCFw69atwtraiYcyJkvVBHfF7ySYMiPwHX03MIMd9TeBKHIwIIsiWBlhY3sb/+FLfwApOJ5/5jyOLBxANug7eSCtEcdRYYCnIJgE2TNoWyglMGdTXuQoaGNguIQ2Almeg/EIIpJY2ejg2t0VbGz38fobb2Cj10N3oKE5R7ffxyDLESVNcBENmZfVLUP63kCU+H2XVN9em6BMH94Md4vqlkv9QOg/l//vQ5tsKmSUZ5sR6qFVJbpJvIfGCZGOmj/sttOqu35H7TSNmzvdD+MwhDGpYKhLAA9qcPcw4LZdHMIY0zDTTugbYPazeEIapQ7nKv3zOVM/Y4X4ZhHFCxRUoihCHMdlR0PLjT5pwB+M+gGQoLg6/TH/gqXEBgBHjx7FmTNnSrbWnTt3ykA5NzeHF154AXme4/bt2+XQnZeyPe7L8xOFZcapVYeQnXVdkoFGnltwzqDzDDNzc1BJhO7WBn7r3/0ubt+5ix/4vu/B/j0z0NqCSYOByiGYKPZ1FLhwQqMuCLg9IgWLXDv/Is0YwBtQSmFtvYs0zzBIU1x69328cekKumkGKRMYxjEwCpxHzsIhThAJOdRt1AWu8BzT79O8ziXPeCg5+N1nOLMBnIKCn1xCWI5swenzHvV6/E5onNDoONfTUVYMu0kQu4Xe7id51M2ERnW0kwi7hojC4wzFjaOOV5xvDoYmpp3QRzwBLRyb1yp7JjPZD2lmv49H8Rkh5AxVrMRuI3w/yzL0ej10u10AQLPZRKPRuCeI+RWaX+FWdUKhlMyZM2fw7LPPIssyrK+vwxiDRqNR/k673cbevXtx5swZbG9vYzAY0AMVnRAvE4x70mJgC+6J6pgySVlmwKyz1WYAokYDaZ6BA4iSJqBzrGxs4erN25jb+yy4tbAmh2EcTEooxqCM66dypcC5hJARjLHo91L0UwXLOG7fvYObt++gP+hjaXUNq2trEFEEywQ0jyFiDisTdLp9NNpz2NjcxFa3ByYiiFhCRBKcu70jY0glorCh8AJTqHRAwSnLsns+I39m48/xQtkeYuGFtg95ng8xIsMBuR8Y/Z8RocV/7BDqqqM+j0pEo5LBqO7jQedAH7QFxbikWLUb9rjAcZMmxntmmgzCWptMZ0IfVeht4biAMYeVyT6bWfUzRvIXwfgCF5L5RALqYrLM2Vqvra2VNN4kSUqJl3IW4rGpfJggXISsEmAEgCzLsLGxAcYY9u3bh3a7ja2tLWxubpZwQ6fTgTEGx44dw3vvvTfEyPPnQYYFueiem5GXCcgWatR5rsC4Ix5YBkTNJrhp4ObyGv7Zr/46/vmv/TpmWk1IzhEXFPJDhw7h6NFjWFldxfLyMvr9PriQYODQBQ3bWgbDrHN+BYMyBorHUEw4IgY4tGFQgwwikuj2ejAM0Np1ZzszuXukSksNOv98V3UV1KUQk5E+vyoVi7BACGVoiMFI3SuRCXzSSB0lmQoWH7Ib1wntJuBP4pD6MBPEJF3NpEF6N3tKoW6cT6d/XGZBD5iguLVoTmdCH8Xu5+CxttH5U7nN/1Jq9Y8wIc8KIdtUQcdxjLiQhyF4LMsydDqdEp6JomioWq6CXXxnTp+gEEqbhMFl3759OHnyJBqNBrIsw/LyMqy16HQ65UKlTz32l2CpsxmCLEo9AwPBvPmG3bHXdhYRBrHkpfcP4xLGaudcGsVQiqHf62JbWbTbbQjlFA/Uehd3e+9BGY1cWViZDHV+nAlYPtyZGM5hOYc2BlZIaGWhrRNF5YzBGoVIMKh0gLm5NiIhEQkJJ+zDhgVPBR8Z8AGg0WjgwIEDQ9bkVd2pD6dRkkiSpCSekJEezZfo8+j1euU80N81CgfpNJPyrwlKYHTNhEk0rPirSC1VqtYhtDUuwU0y8xkFy9Wd+zqbBX+eVvXaqdsclfDCz25UYgqT0yQQ4YMmlCpCQpWyR1WCtW6Pu2XtRyN+T5NQcZzcf2Qxywd/Lof6y0bw75Bx4whjTNBFHEVRefFTIBkMBhgMBlBKlfBcncz/brfZqzDuKIrQarUwOztbzjJWV1fRbDaR53lJgqC9l1F0Vvc6CJ7QpSGeby630/2zoc7JzXUkwA0MDAy3YHETqdYwgxzNZhNxEqNnAZEXgpw8Kky5vODnme/t3GTkIYRCEFU5RQWzQ1/O8xycWWfVUNGpjFru9P9OiSIMbKN2fvzPkWBZ+n1i1eV5PtT1jqOIh59znWL2pA6hVZDfpJX2bqRuxiWlSYLzJEmt7nl9YkeY1HwdPv9n4yjeH8QxSRe3y5mVsNa2MYXjPhrHqYPHWkar05kefF9u1Q/xOH4miuL9PpRGwcrfmKf5D1GmqbMZZcEQ3mB1StnhRUkBLc9zWGvRbDZhrcXMzAzm5+fR6/XKqi5JEqRpWgZIkggaJQm0W6kgvyKlG4xgKFqYJWjKV4TwFy7D/x7l9RKqHfT7/bIoqFryHcUCCytNP8H4uyg0rwsfPwwo1LHQ+6R/TzBtSFqoq4RDOnFoke1/v6qoqVs8rWNeVqkNTNLNTOJltRvJoFHX1250Euvet49A1HWOdd3lqJ9/GIdHsuAAmtbaaSf0xCegA0cXtM5eTHX6Vwxnf17EjcOM84Y/K6D5DwWjLMvQ7XZLif9ms1nuAI0SGw3p2GE1O+qG8xPK1tYWDh06VC5VtlotRFGE+fn5shK/fPlySRGfn58fqgirbqSQNh4GoaoBuf+efBFWEv9USqHVapXwJXUck5izhQoC4VeapuVCaZ299qQzi6r3XiedVHX+iERANHr6e1Z4RlV1YHXJkq45H4YbBd+EzK8wqY7rIib53VEJ6kEEUEf9mzqrhyqYbpKDishQkaLOMPBhwXCTwnT3wdwTFrZlPyIW39+QSejMwvGG0eqEMul3ZVb/hI3kx6SM9vkVvg+v0QXc7/dL1pkQwsFOBa03nCNUJSG/+hy38R4+jhACm5ubuHr1Kg4dOoS5uTk0Gg3MzMzAWosjR46g0+ng5Zdfxte+9jV0u120Wq3ytY7aQaqrpMPOZdQN43eBlADpcWlG5m+wV8nQhEwmGu6HSYhmXaH30iRaaqMqdj8gTyKRI4QomW+k50fdk/86q7qvOoiNNP98j6NJO4Y6w7tRAXCS361LOLtVDR83O6rq7KrmJFVFx7jnps+k6rFGzbxGwZMfhJL2KLsR779ZoSCeTJPQkwm/HdA6fz632Y+lRn+3iOLjQoiGj/1LKUt4jYJBv99Hp9Mp5XAajcZQ4A0DWN2NUiXHUndR+79HigivvfYa5ubmcOrUqfLGajQauHPnDl577TW88cYb6Pf7ZZcQx3Ht7gm9Lqq+Q7inahAevmZPWLK8iagzpP2bdrs95MMTqkuEmmphwqHn8wf/VBzcr3FZ1Rxh1AC5LkCFydtXyfChyHGdg3/tkThnOM+o6oyqlBwm6XB2Y2swyayj7r1N6oFVlYD89+Yn7bDwqJNPqjqH/pxuEuvxUeejTul81B7TQ9xXSoBpEnqijtMLJ0Qhu/PZHPonLecvijhZCCtzIiHQwDnP81LckggISZIMMeD8myL83jjnybquKazQad5w9+5dvP7668iyDEIIpGmKwWCAO3fu4O7du+j1ekMMLFJtGDUcJdUAYvz5QquhuGrVzeg/PiU+VmjBKaWQpukQtT28uauSmv8afGaYzyykz2jULGAcFBTOXEbZKYSPTVp3dA7pPfd6vUqx2klmJFUsvFEGh3WfaUhueED4p/IcjJLhmQSum4RO7pNERs246q6pEKIMl4pHzdN2Y58+SaJ5WPJLzHl5xfiIGNt9QySh0wePN/Osf04x/VMK5gtMyFNciGYVjBYqHOR5Xkr7SynhC5VStxFCGlULkeMqyVFwEf0OkQ6Wl5fRarXK+Yi1FisrK1hfXy/9bupgqqpAVGVXTTR0vyoNVQl8CCusiGlfKsuysnvxE30YKMfJ+ftyNv6czhf1nATyGRVQfMUCv5r2z09IraZO06df05JwlQFeeK3UBVZ/V6hudrFblYNJ9oImsfWedIg/Do4LE0Ed0aJK8mg38FZ4Xkd1Qrud5+yGCTjp98fFi0KgNwLYNAk9EfOfg0fns6z/8Qz539CMfT5KGkf8i8+Hh8hXhoJev98fsniO47iE6vwbsKpTqKqMCLIiCq9f+Y5KQP5NGEURtre38dprr92TRGj+EA7J/QDrw1v+hn+j0RhSCTDGYG1trfw5zb7C1+bDJGF1miRJCWXScxB5Ijz/VTMN3+q61+uVpId2u10+Tp0KwaibOzy3Yafl+/nQZ+8nTn/J2FdKyPMcgNsd85MkdWx+Re6/V/+xKXl3Op2yaxwFG4X2EnXwb9Xv1fkbjesKdgtNVTEAq673UGE8fBx6D81mc0jmiHbifFjYF5j1DQvp8wqvW3qsSYguo8gqdTtOdXO0qnMzSnKI3oeQIuKGzR/bsyBvbC6paRJ6XBPQgSOLeT74thTq51kc/7lIiL1+EPGTj09GyPMcW1tb6PV65YVNNGxf5LLOjrsOXw+Nz0LpnlFeLn5F7UM2fuAM7QD85BPOvPwbhmA7IhMQ3LW4uAgA2NzcnHhOEgbGOI5L6nae5yWrze9ywhvOD5z+bhDBoZQQd1vF1llL0zkkiR2fDEGdJXU6PhNQCFGeM1LPWFtbQ7vdLq8jrTUajUYpTkpMwaquyO+ewq7MLxp2O0yv6jon2TOq66DqZj/jiAaTQHdhIK7693WFR1XCGEVdrztP466tce/lYUNwNVdzbGHmihg+TUKP23F28YTUKjuZ6fR7Uqi/zuL4OcZ5M+x8/KBMwabf7w9RsGk+RIGZklAVhFJX4dVVO+FAfJyQqX+j+NCCP4D1Oyy/Q/KJA8Q6S9MUeZ6X8BFBXSTKunfv3qFB7jh4MQykYUVJ3SWpT1AHUgXz+QHHTw5xHJdB/UFveB/iaTabZYKhc8I5x/b2diluGlbntCBMHdpgMMDc3Bx+4Ad+AK+88koJkfpVvN/11OnC0fVGPlR0nnyZoDC5hEXRuOBZFejDPaLwmq7brxmnbTfutYyCt6pg7fB6qSIyVCkx+J2Wv4MVLrCO6u6rXu+kkNqDzOLuOS+cSRjMA4gADKZJ6HHqfhaON1SWXshZ/tM5sz/CouQkY0zSh+nL2PhMOGIlbW9vo9frlXs4PlW7SgBzkqXTUZBEVfVXV91WyZv4FzZ1DeHMxE8ApPBATLPQQI2CK6lyhyZuVXDPKGkcqvybzSa63a7Tj/O6saq5R6hYTa/Xp2ZPgsdP0ilxztFut3Hq1CkcP34cMzMzGAwG6PV6UErha1/7GpaXl0sINhxs0+vM8xytVgs/+7M/C6UUnn32WVy9erWEIkNW4KiZC12TtJwczvKqoLgHHXY/DirTdYkuPKgYrLJnqAr6Pvrhe0BVdU3jPJVGzeEmLSLH3S8TzqIkY3buoxDDP1JJ6MzB40mW9j+WQ/2ckfwHRJQcDeEvP4EQ0w3AkA0DVeq+oVmdCkLVwHrSimaUWkDdJn0V3ZpuREqwPmGCICGyAu/3++Xv0nsMvWuyLCuDri9FdL+DVUpEcRyXiZAgzhAqqkq6aZoOwYs+LXwcDDPqMMZgfn4e58+fx969e8vkvW/fPuzZswdRFKHf7+Pll18uTe/C68m3gPj4xz+OVquFbrcLKSVmZmbKWVuoV0Y7RnXFSAiZVhUAVQXEpAuok0B6u01go2C3UcF9lIlfHdxL88Ysyya2Qhhnrz7J9f0gJIb76X7qd/i4BNOz+AioJnxkktDpA8caWdp/IbXZ37SR+EEho0X/Jg2TCAVFzjl6vR56vV651xLuCYVJbBStehQdNZSgqdp4H1XN+QnIfx5f2YE6h16vV8JtlFj9StuHI8LXTzc5dUH+HGxSVlBIUSZ3WYI8O51OqahQt9tCwYE6sypx2Ekqx6rXSkSJY8eO4eTJk+Vr8eE5zjnOnTuHtbU1XL58uexMfAt1IQQajQbOnz9fejkJIbC+vo47d+4M2Tj4RIYqmMknlITdYRXjsmrvLEzqdSrgVfOoUQK6k1TrddBcnavrJMmw7qDkTpBlFUQWJpoqCaiqQjCcOYXX4yQdT9252u0KQS0cx5iwwB477YQej+PU/qONLO2/mCH/OSP5D0RxsugHVPrwKSBSkuGcI01TdDqdezoE366has6xG62sEEILZXTq8PEq6M2nkodBhZh8WZaVCSh07qyrsv3gkyQJ9uzZU7IEfQhzN1WeLwLqC34SSYHmbqMSEIAhwgQVB3WV86j/9gODUgr79u3D2bNnEccx9u/fj9OnT2N1dRVXrlzBYDAo3/e5c+ewsrKC1dXVIXZVo9HAxsYGTp06hZdeeqmkzKdpinfeeQfr6+tD7D+fzu/DnGFw8/et6hiNVX8fpc83KmmMmyWNCpIPMucY1w2NUmkg+n/V+ahjoFXZvFcpiO9m3jOKBfewZkKV8zE3Ypiz1sTTJPThJ6A4zwYfy5D/TcTR90dRtOjffP4NSLCSv9G/vb1d7tpIKUsacVX3U3fDTuJOWXXR+/+GhtyjdkJ8CjYFMko4RGH2b0J6H1WsKj8x+XMXOgf+vpE/gxkX4Kuq3pDZRB0RdWm+02xYyfoq5T5N/H5val/V4dChQzh06FBZfJAtR7/fL6+JPM/RaDTK10wJiHOOzc1NzM3NlZ3U8vIyjDHlMrFPbQ8Lj0kCDunuUYfuL1z6EO2oJegqNYW6Dmg3xIZJupe6RDKppfco9hsViXU/9+d1YWKqmguN222qS0APQ19uN7uE3n8LY+2sMXaahD7sQ+XZmYFJf5o34u8RUbRY18KG2/9pmmJ7exvdbheMsZJxFdK3q4gIVTfuJNULBQ+ClJRSZYCn3ZJwM9zvQijxaK3LTmdubg779u3D9vZ2GUD9uYNPAffhsarZFM0xms3mEBNr1O5T3U1ahcX7v+8rg1d1mXQOut3u0A6X/5rrgnoIcYZsMmMMDh48iKNHjyLLsnJWtrq6io2NDaRpWnYfZKPu76HQLGJxcRHf8R3fgcXFRWxvb5dMvrfffhvb29tD/k7+7C2UmqnSRaMkRJ850bvD3aQ6LTX/8H1zqs6J/9yTzJOqguL9kiTqZh6jCg16nT5VP3ysUCHBP+e+rNJuF23HzYsmMS6s67ZGMRb9wrp47dxY27bWNqZJ6MPsgvYd2Zuq/uetFN/PZXTUZyGF3RB1QcYYdLvdcgZUJVYaCmNOIjo6brkt3H2hAEyJodVqjbzAlVKldQQFQQD42Mc+hk984hPodru4dOkSXn31Vayurg4lvTBAhBd7lmVoNBqlIrcf6Cdl7ew28JDsDkkGEfxFQd8/D/S7IQQ5KfstHO7T+SBaNT2/b6XuLyT7wczXq/v85z+PkydPltdSv9/H0tIS0jR94GG2T1Agphwloip175DCHy6n+guaVR3UKOhykop/FPlglDJIFZEhfP1Vr9G/hug+Ggfx0WfvJ+OHzQrczeM9CCuRM8Y10LJAa5qEPtwu6PhAZz8oW81joUBmGIjoe2QGR4wrCm70VVfRjTJOGzeQrYJQSNONGFQhTk1QENGoQ303XxV4fn6+3OmhjogSXRiMqvZ3CLqjTiOc5TzsBORr9BH7jYRhfYiQzgHNgnYzg6ur2ikp9Xo9bG1tYX5+fojQQYnOD3CkXkALp1prnD17FmfPni2p3MYYrK6u4pVXXin1++q66HGdm59MKBHR8mvVEnJYbNRJ34RfVYkqfO66Gc44yCyEZ+vU2OtIC6PgPn8+Sp9RFcOyinxRFR/GwYd1heXDhOCqOuQJBkQNMDSnSehDOk7uO8KzLD2pYM9EnDerqvdQEZsqXtrdoM7HD351gqSjYLZJcG7qgHy4gMzxiKob6mTRAN+3kPaXThljWF9fx+rqKg4ePIjFxUVcuHABN27cwO3bt8ubtC5I03udnZ0dgrqqYIEHqfaqZmKhcgN9NjSzoyE/KQ7UmdeNq0SrxC+ttdjc3MTq6ipOnjxZwmYEyfpBOoqici5Fj6e1xuc+9zkwxsqCJk1TvPrqq7h+/XqZ0KsC425nVzT/oK4xFJmt6oCqbCB8071Jdo2q/KXqGHpVlPFxndK462VSWK6O5VnFPvV3tar2vR40sdyva/K4e6oOeuaCRwBaJw4c4ddWbplpEnrUXZBSjUE2OG2EnaUFzfCD8xluWusShiM9MKqwfcpyHRRXp7NVxcypqvSoiqZAQclhMBig0+kMQYdhNeTfbDS/ok7n8uXLWFxcxKc+9Sm0Wi0cPnwYzz33HDqdDnq9HrIsG0ow/nug995oNO4JSFUb/Q8DlgsrY/ociGRB55+6FWIrEsliVLIZd9CmPCWPtbU1dLtd7N27t6Rk+/MTay22trZw+/btsliw1uITn/gEjh07hmvXrpWqCktLS3jvvffKc+o/zqSJaNRwnhQmfDuCOup5lb2Dz8wLi52qLj/8fX92WDXnG6U8Pioh+cSZUZ1PeG/Tnz5ppkr6qSqg+/OiUWod4wrPUX9/kG6oLslXzABjbXXLWkgA2TQJPfIkpEU/6+/XksdsMCirZT8B0YdGbKdOp1MqCiRJUi5rhrOCqgsq3KMZdYFW4dy+W6bfEfkq0aF8v0+S8AUZrbXl0LrX6+GVV17B3NwcnnnmGczPz+Pbvu3b0O128frrr5ddX5ic4zgu33+du6k/P3gYGHl4E1Og86EvophTsA0TkL+sOslN73dBoRLz0tIS3njjDVy4cAGHDh0q50BE/FhdXcW7776Lq1evYnt7G81mExcuXMDnPvc53LlzB4wx9Pt93LlzB5cuXRqizldJRI2y9K6jDfuv2SdJVFGLq0zt6qR66ha46wgL4XVQtzdXR9ipW2vw5aZG3V9VcJx//4QJNRT+rSqqqmwdRjENJ50P76ZTr1MhqeqIK55AGq33wDmsTpPQoz6M1lEOM6eVia1HMKCgTd0NzYB6vR601kPJJwzydSy4unnKbvTUqNrzg75fhfkUYD9I+M9JcyD6t0IItNttLC8v44033sCePXtw7tw5HD16FB//+Mdx8+bNUjHBH3QTBduv/ENJmpAO/KBJqO58AhhKMmSfTgrWVFyMgtnGXivBQJ4Cer/fx+XLlzEYDHDw4EEkSYLZ2VlorbG8vIylpSWsra2h1+thYWEBzz33HD75yU9CSomtrS10Oh1cuXIFly9fxs2bN4c+sxAavp9OMkxMdI0TfBmK39Z1AGGArptz1i3Q1u3SVCWicUKnozqC0LJhVALzixe/MKk7f2EC3Y0ixLjv3e/C7W664prXEGut5601T/Rs/8lNQtZGBk7Aj+YnBDH51ZCPAYfsN5/I4N/oo3YaduNP498IPrzhB46wovcDWBWM4GPvFJyllFhfX8e1a9ewd+9e7NmzBydOnMCePXuwuro6pAjt7wD5bEIfsvLb/jAphYFoXEdSVyWHla8PhSqlSmiuSqzyfpw/w6Evnb80TfHuu+/i3XffhZQSx48fBwAsLS2V1GitNZ555hm88MILmJ+fx/Xr16GUwq1bt8oE5C9DhzJPdTOL8M+wI6rqHCnw+tbnoxLBuCBXN/sZN9OZRLl7XEEy6rWOIxn410yr1cL29nbtufW7Lvp3tBNHcWHSVYu6e3zSBDTO56ruHgnvH2stGGeRZdhnn3Dpnif2xVvYJoB9UgjGvIXLkMZKg9xQrDQMcOOqo91Sg8Oqra7y9H1s/GBTNUugIES2CwTLtdttrK+v491338WePXvQbrcxPz+PT3ziE9ja2sLdu3fL7om6QKK1hnMgStS+Ed2oG+V+Tb2qOiR6bkqajUbjnj2pUQZx45JRnT0GPZ9SCktLSyWES+dmYWEBzzzzDA4ePIjV1dVyp+jtt9/G3bt3h1S2fbuHUYyy0BxvVJIICS7hebofEc06EkHYOYyzKanqOCcp0MYVbnUJu2qW1Gg0sLm5Wdt5TuIE+zC6l/uZA+3m39x7zbAIsPPTJPThpaGmBGaiJBH0QRGWPxgMkCRJGbB9IoKvMB2yhOpujFE34qgLvW6gOwpGCivpcHmT5lnE2IrjuNR5u337NtI0RZIk+K7v+i58+7d/O/I8x9e+9jVsb29XUmXdfE0NbZ/TrkxIK/dvCJ8SvxvILgyqobafv2gb6sTtFrbw/ZKqAjXBkb6/D4mPEn18a2sLP/7jP44jR45gY2MDKysr6HQ6+OpXv4orV64MLZX6ECvNHuvmEHXstnHq5PT6iYhDsJyvDvAgNhdVCahqt6iK/j3K3qQuAI+Ctuuuq5AM5LNGq4rEumvO74weBjvuQWG2OpJDiMR414nQ1s5N4bgPKwVZ2xZSzkZRJEM7g263W84afFdPP9BRwKhjwu1mADkKO/eZSVVBt+p5wjlVeKMSBEEwpBACzWYT29vbWF5exuXLl3H+/HlEUYROpzM0S6hiSdFjSynL/alGo1FSpquS5Dj14fuZGfkDfHrNVdXtpJ/BKEtzH5Lz52x+kMvzHJ/97Gfx3HPPYWtrC8vLy8iyDK+88gouXbpUvkbf7p0O30217hyNUkUfl4T8zyVUABgnAVOlwF3n6DlKuHfU/XK/1PRxxV3YqfmGlNTdTzJbq5OgepDXfL//dpzKQp3xoTFGWtgZa59s6Z4neCak9zDOZ0O2D8FyW1tbZSXqExZ8h8tJdNEmTUDjBplVEFxoLVx1I1fRSf1ZF23nU2CSUuLKlSv4wz/8QzQaDVy6dAmbm5slPTmkOdN7TtO0hHjov31ZIQrWdSoM91sFhkNjf97lyyxN4jUziRp5+Dn5S78ECdJrOH36ND7/+c8jz3Osra0hz/OSCUcaeH43RftN9FnRdTau66hKROOG334SpaTiO8KOUhwYNYvwr6W6uVGVDuGohDtKfWHUPTeK4h1KIIX+S3Xdt1/sVJ2nD/MY1RXWdJcCQNtaE02T0IeRhIyZZ5K3wouOgiYNlSnAE3RFNy2xxigRVWHJo9QT6oaSdcPXOojOD35Vz+EPYP2DZkh+cojjuITprl+/jizLSidTHzrzAxWdC8YYsixDu91Gq9UqYaaVlZUhyMqHjfwA+CCJqOpchfJJk3Zd4wQpw8NfFKZ/F0URFhYW8JnPfAaNRgOrq6vI8xwrKyt45513hroegoLCLozO6ThIkkgYoep11WJp1aworOxDp91xRdKouU7dML7uMxyVXOoSahV1vW5Voqrj8pMQvf46RfaQeRp2j/dTcD5qM8CgQBUWaJonXD/uiUxCi+39Sae3dYTzqFF1Ifg7QnTBkUxOKBlDQaguCYzriOr2g6rgpvDmCQPJqBkRJYsQEiMIbTAYlDdiFEXloirBSkRioArXT860f9Rut3HgwAEcP368rPJfe+21Ul8tZOWFskAPCmGEcixVxcHDSkChsjfBtMSQu3DhAs6fP19SsVdWVnDlyhXcvHmzvJZ8eJR056iDq0rOIWWY9APpGqyixVcpH/iQmh9YSdx0UiHQUeKdVXs74+jXo9CEUdfJ/dDYw+6KZsBVthjhuQtp7eHX/ez/PAgUNy5hV3mRlT/nrAVH0pomoUc8EIotzKIQIvbnLbRV7tv/UsVKpAWlVCnNT+KdVTpau5Gsn2Q+4fsShcPnUYSIsPOpY9sR9EOdjA9NkCUAPY5PPKAkpJTCSy+9hJMnT6LdbiPPc8zMzODkyZP4kz/5E9y5c6cURqVze79Q3CjKe2iFPQ4erTIwm/TzCT2dOOeYn5/Ht3zLt+CTn/xk+Z7X19fx8ssv4+bNmyXb0idNUCIaxdirsi7PsqxM5JR0/cGzr4xQBY+FpBB/3aDKr2qUrfi44oBgxzp7+7pFVz+x1pEX6pLhJJYP9H1aavaJNVWdp//4PqGjzjn40Ye28S6xw++HxQCmndCH8EHFYGwfABni1b4AZThDoWBNdgdJkgzZBPt7Rv5NRrBe2PWMYtaFWG7d706CifustpC5Rl0MqWBTwgkTFQUxCqJUhZNG2+c//3l8+tOfxoEDB2Ctxd27d5FlGWZmZnDixAn0+30sLy8P2ROMg+Gq7AqqqlgqFvz5FgWUqvMyytkzfJ4q9YAqjyMqXj7zmc/g1KlTeO+99zAYDLC8vIyvfvWruHr1KpRSSJJkyPq8Smsw3J8KkyQVAlQ4EM3e/4zpXPj0cX9e43eN/uOHMF6Vvhv9XhVMXNVJVMHTdQuxfmdZda7H7QjtZv8mvKdICJju17Cjo9fod6ohg3I3zql1gqy7KVKrqOLhGsI9+0F+McoQWdjk5IFF9v7KXTtNQo8uC0kAs8y5C97TvfiLqP4F5gdPgqoIovI7jjCA+bDQOL2scdh5VRAeBeeN6p4I0iEVBNKAoy4oDAb+DUc3IDmHfvzjH8fCwkLpqEodQKfTwdzcHGZnZ7Fnz57S34dmHpNUbuN+Ru/Zh0ZHKZqP6jCqEnoII4aafICz8/7Wb/1WnDlzBhsbG+j1elhZWcGf/MmflFRsosIThXvS5cyqLojkiWZmZoauQUrKpGtI3ToZ24XvoWqGEhY+xpg+AM4YixhjPEzIo8wKq+ZFIcOzao9nUphuXNCfRJ2E/ptce0NI00/+ofqG33nWvfdRDq+PwRFZaxJrrQCgpknoUeUg2AhAi3F3Q1XJeoRwTojfk5wPDfTphqcA7lt71wXOSVSdR1WOk4ofVlGN6aai109MwFARIGR/hVAU5xzHjh0r6dwETaytrZW7RVEUYc+ePVhcXMQ777wzdC4flKbtz6cI7qFz7weMSayW65JbaK3ud5Z5nkMIgaeffhovvPBC2ZFtbGzg61//Ot56660SwvVnVXWw6bguze9sCCqm/bU0Tctr16fLU5FBnatfwdct8nqw3DaA6wC2rbUz1tojANqMsfh+5jJ1UOAkxdekCeh+FzpJgd03JaQCkq4t/9oNnVknKSoek8QzFMOttU1gmoQedRaSjLMEYLwuKdRtyPsyPuTRQwE9SZIyMBA9ObxQQ+md+x1KPgyzOH+fpqp1rwqCVRbfBw4cQK/Xw9LSUpm4tra2hqrLJEnKQEyJb9K50CRVNs2mKCBPuvlf91n7QcOHL6ga9iV2Dhw4gGeeeQatVgvr6+u4cuUKrl27hvfeew/GGMzMzJRBLEmSoaXacXTicPZBXZBSCs1ms1TvDhcnsywrz33V5+kXEVW+T2US0rrHgFc58DKAHMBZBXxaa32WMTbHOZeTFFJ1s7swGT7INV1nilf3s/Bzpnu33W6j0+mUcGdVXCDldh8RqILcxiWjR82OC18X51zC2tlCNSGdJqFHloPArIUAwOoGpFVmVv7F5icX37WSHE5J0dkX+6xj0TzMim5S+In+Tt41YXfjL1yOsxPYt29fyYAjBp4PXdI+ElXmROqYZM9iEvq2L68U0rJ3m+BGbeX7VHUqPIh8cfToUVhrsbGxgffffx+vv/56qbxB79Oft4yCC+s6V0qCfkKjZE6PPxgMMDs7izRN0e/3h7rN0CtoEpiTAUoC78yK5u8ILpa1MUlX934rA75grP1+rfUBzvkM55xNAo+Nmo9MkoTG3TOjutlxmnbUqTabzfJ69q3Q6XokSFVKiSzLygKojmDxsO/fh2mPwhiTsHYW1nI8oceTLPdgwyqzbkZDNy8N1f3KiSohrXWprkDDZ9+P3t8xGrWZPglt9WFVQX4wDA3zQu+ROgMvY0xprU0UX4Kf/Jsmz/MyIFNApQXBSZwqRyUN6g78DmU3/jvjpHvCIE4Fx/79+/Gt3/qt+OQnP4k8z/H+++/jj/7oj/Dqq68OMaa01uXuFF0fVTOHuuf3ITiapZGYLCle0HV2/PhxfOxjH8PS0hLeeustdDodpGlafqY+m9Of8dV1YIwxJi1WkiS+eau3uQ4Ahxp7budKvd1V3T8bAD9pjHnOGjMrpJyZxIp7HJkmJChMOtupu8bHFXdh0qIVDCqaqmbCfsFD5/6RBq+KQvZ+4gTjXFijZoqZ0DQJPcLDAFa7PyGqLsaq/ZyadraEs5RS6PV6Q5Uv2U/7ezYPAjOMS1qTwBS+MoTvMeRDW35i8N04qzbHL168iAsXLpRQVahB5ltj+ArcPizzIBAjCc/Srsck1WidFM+ortFP3AcOHMCLL76Ic+fOYXt7u2T/LS0t3TND9LXJfJPEST7bMAkR5EhJnkgOg8EA+/fvL2nyt2/fxp49e/DWW2/hvffeG9r58gkVo4qe4meCgYMLXvrN3Bls5gCuH2rO/8pgMHilawd/MQd+SCl1inO+h3OeTHodVxEcdtPJViWyUX5dIfOzLsG1Wq1SiJYKNJ8m7iumhMoWdRp0j+khADSnSejRHxoWBPgOqQ6MMtsK7Y/9ISsNnMnhk+YgrVYLzWazZCj5c6NxN9Nug/IoxYWqgOMP8/0FUn8BkmDHkCbuw0mDwQB79+4tteJarVZZaWdZhtu3b+PatWu4devWPd2Vr5F2X9VE8R784f9ug9eoBOV3i7Tf1G638eKLL+LZZ59FlmXodDq4efMmXnnlFSwtLQ2JYpI8DyVJcmX1u8K61+InK//nBBn5nczp06fx7LPPYmFhARsbG2g2mzh27Fj5fDdv3iwfh+jbk/gpMcaktWaGVXxAd/obW8dmD7ya5I1bvUH/q32kX1DGfN4Ys0DJqIpBV0cvnjT57JZVOUphIYTe6XvUuWqtMRgMhhKYrxhS9b1JlcA/KHhulwUus9Y2pnDch9AJMca0dXdCrddNWC35F5iPtVcZghFERBAd/T7NTHydtaqN8vvFleuWL0PJHILDer0erLWYnZ0dgh3pBvM14Ki7oSRK73l9fR1LS0vYt2/fkPozdVs3btzA3bt30e/3h/aExnUh4d9DxWL6IisEXzl7nPin/5hVqgL+Z0xQHwDMzc3h+PHjOHjwIAaDAbrdLlZXV3HlyhXcuXNnKBlScvc7RP+zHxUsfTUOIhqETEzqihhjaLfb2Lt3L+I4xubmZtlxtttttNttZFlWfi6jglj431xwwWD3+oiBf9zYXrEAlo7OHvyDRpZd7KTd306hfsAY8x3GmEXB+SzjPK7qSELoz+82qmSHQsbqKJhv1D5O3U5WuNwdRRHa7TYAlOffh5x9Sxe6R6jQGOesOqpTGwfPV523cTO3OuUMay0DEFlgmoQe6cGYBaAtYNkEuLzf8YwyFaMAQ9UmQV00wKaLm/x2KKD7w/8HwXdHVfRVAqd+UqS9Ehq4+nsR9F6qZkVCiFJ5+/nnn0ez2cTm5mbZNdy4cQNLS0vodrtDw9sqK+lJO5UQLqsSRR1Fya5aYq3aFyKYpdlslp3M4uIizp49i7m5OeR5jvX1dbz99tt47733kOd5SfLwSQw+PDiJdphPofdhU4IziehCn1Or1cKePXuGKvNer1fONYig4BNHqtxm6+AaY0wbwEiRy5vbyymA60dmDq5lWfb2IOv/Zg/ZF7Qx38GMOSCk2McYl1XLp1Xmc3UK3VXXTNU5HSd/NaqL8BmsBHsKIUopK0rwPlU/nBvVzZvqCoD7vd/HxYoJOksGWAlr2YfB1PsGnwnBALC7CXrhjRNaG/hdjN8NULCamZkpJXGoqqUEEA4260zD7idYhxU/VZk0+9na2sL29jZarVb5RbMGIQRmZmZgjEG/3y+XJP3kJaXE66+/jna7jWaziTRN0W638e677+LmzZslpBTq8Y2r4MYZ2VGC9830fIYSdRLjzpn/eYYVI0FrMzMzOH36NI4fP44DBw6g2+3izp07ZQLa2toaglqr9AdHBaOqGZRPCyfmFlXaNCNqNBp49tlncf78ecRxjLt376LZbMJai06ng/feew/vvvtu2fnSXGhcp+iPrhlnLWsnq5RvdZa7AN49MrNwp5Glb/az/m8NkP2oUvrbBDOLXMq9Vdf5uI7A//1xc9FJRW7HQXe+HQh1QN1utxQzDj2xfBJD2I3vljn4IPf6LityAOAWT+7xJLPj9LhPs8qDxK9ofTFPukFoiE8VK7XuaZpic3MTAMoZkVIKs7Oz9wh57vYiGzfXqAu8dCNRYOp2u9je3i6D3ezsLJrNZhncW61W+Z57vV45A+Kco9vt4g/+4A/KBEfBOPTK8WGo3bzuuvft22qM04qr6naqpGt8Snq73ca+ffuwuLiIkydPlvTy1dVVvPrqq3j//ffLHTHfv8if+1WxMEd1vSFJhAqWZrM5BFNR10o0+5mZGayurqLb7SJNU6ysrGBtbW2IGUcd1S7Uy7kxJqqD4+qT0VIPwLXD7YMrSZpeTFX/xb7Nf0bl+fNCiINcytmwewg75BAmryMe3K/T6LjZqQ8NNhqNMtHQzJTOaxzHJflo3NrBbhPRB0luYIzBAgyuwGDTJPRo8TgHxwWwTB1MM85wrm7g6rPCKAisr6+Xuxxaa2xsbJSabeE+ziRLb5PCcWEQpselLixUAs+yDKurq0NzCAp0tPtEAZA6I6oWaU7R6/UwNzc3ZJrmw4Pj1L9H7XsQXBXuB91PovbnZL4VQhzHOHDgAJ566ikcPXq0DEBf/OIX8fLLL5c7YX7CCZUa6kz1xiViKmiIUk07QQTpEmHi05/+NI4dOwZjDFZWVkr4aGNjA7//+7+Pzc3N8hwRndufR44LUowxxjiX1t5fkLrdXe4BuHSoffBukqZvdFXnc6nWP2m0PikieZBz0aizDfc76LBIq1oA3223MUrgNJyhSinL+dDW1lZJ4KHPhhiaNK/bTTe2myJzUqmn3TZDT2wGenJnQrAEx9VVppPKrfsfut+a+2rTNLwk35c8z7GxsVGqcRNbybcfGNcRTMoOCokTVcN9SpT+cp5vLZ2mKbIsQ6/Xw/b2dpmAqDqXUmJubg79fr90oFVKlQoC7Xb7HhZeHSQyyqysahbkq56HwSMkfFTtZ1UROGggvXfvXpw7dw579+4toZi33noLFy9eLLsS/5rwGXG7kQiqKmLovdF1QUUKDcgBlIuyzWYT6+vryPO8pGtvbGyUj02kCPps/CH7BEGLwULaB2RP3ekubwF4c6Gx70466H8lRfoDWa7+IpM4JaLoIADmQ49V59CHcauEZXfjYlyVzOhndG7Cn0kpS7iZZpw+EYVef51F+sM47gclGaWNOIzKTZPQozwsnE6SnfSDrCIlhImpSmKefpfUE5IkKWcrdLFSN0EsryoK98OyDQ7nIP77IniHqm163eEFTZ0PUdEpic3Ozpa0bKraZ2dnhxQNKDkTdFXF2hk3wPUDUah9R4/pB99JukRfK29mZgaHDh3CoUOHsLi4CCklbt26hddffx3Xr18vmVBERPCZg/71spuAEe6xUDFAS6nUGdD7bzQaOHv2LBqNRvl6hBDo9/vY3NzExYsXS+YjdVX0WfuSM+O6BMYYwMDvtxMKj6XB2tqxuUMbSZZdT9P+Fweq/1dypb5dxPExxvlsKJobzoGqOqJxtg6TLDyHv+93xVUqJ/58NSTt7MZb6GHCbSHMPKEKhQWYKdChaRJ6dI0QDMAUYM39wFtVWH94+EoElFwIlpqZmcFgMMBgMCi7Dl8exK/46E8fKrvfmVEowBnaNPhWDdRdEBRHUBRtkVNA8CvXwWBQBk1/x8afQRBDy5+j+eSO3UCPoUV11aynqiKsSsj0Oolptri4iKNHj6LVauHWrVu4fv06Ll68iDRNyx0fSkChF9AkVuL3BPqgw6NZl092oHMdxzHm5+dx/vx5CCGwvb0NKWVJxNjY2MDVq1eHkjLN9XxLh11eQw8tSN3YumMALB2ZWViPBvGNvur+7iDLfpYzdkEm8SIXsk2vke6LEMKt2uOru34mDfShtFG49xMueNP1S1A0FUIh9DxOfPhDrsctgNyNh6ZJ6JGeeaN1zq078aNM4mzFHlGdaV2VC2SVfwtjrGQw0a7JwsICAJSJiaATonT75IUq3/hQgqUu4IamZb6Ei8/o8t8PQUE+6cJnAimlsLW1haNHj6Lb7WJ5eblkAtJ7pVmJlHJIwsZPTPQaqEuqqyh9e3WfDBDO6uic+VbZvs5amqZlojXGoNls4tlnn8Xp06cxMzMDxhhu3ryJr3zlK6UYqZ94KFn7u2N+gL8fzN/v8Ig2758LIQTm5+fx0ksv4eDBg6VHE3WmBMXR7krITAxtOUaZ/BWvw3Jj7QdB373VWcoBvH+4dWAlGfS/3jHdv9AfpH85Fupk0mwe4FJG9DmGNiI+Bd638Ki6Fuoo01VkoFBY1i/gqNAiQg6pUNB+ECED9Lg+CWTcEvq4nZ86VCCc8Vap3dfNvgtigmWMpYwxM01Cj7YXMozxtJgLPTAuOyro+N0GBU+6iXyMfnV1taRH93q9MvgT8yacedRV+OOSkB98fJjDZx5VeQnRzUauqSSRQ3pmAPD5z38e169fx5tvvlmSLqSU6HQ6ZQIiyRmiC9Ngl+zAqfr1E5Ov3EBJi2w0Go1GrWo2nW+CziiBUiCZm5srz//8/DxeeOEFHD16FPv370en08HS0hJeffVVXLt2rXSKpS6FOkRf0eBBq1tiUQIo/Z38a4uKgP379+P48ePodrtDC8VKKXz1q1/FG2+8UXZGowbku0gsZlLo+n6O272VLoB3FpL5u2na/6OuTn9yu9P5i7EQhxrt9n5/OdqXMAqJJHQO/c62CqrzNeCqdpFGaekRZO17CxE8HcJ3dQlklC36B9vzVMpSGQA9xpiaJqFHmYIYNGPow30A91Cww2qhLsjU4c/+UNyvtvwbJdyXoWBObLnBYFAGUarUq9wRq6yYq/Dhuqq76r35CSjUyiLlYH+HQkqJJEkwPz+Ps2fP4qWXXsLFixfxa7/2a/eoD6dpOiR46jMIfWVyznnZLfpadBSA/H/r/6wK6qBEQeeZBsxSSvT7fRw/fhzPPPMMjh8/jna7jbt37+L999/H+++/j8uXLw8xoDjnaLfbZTIMi4O64FJn8hbOGej1UVKmx+z3+5ifn8dTTz2Fc+fOAQC63W6p+CyEwLVr1/Dmm28OdUEPTdX5EQTKpXRj49jMwT9tZPm1Trb1bwZa/83O1ta3ySg6HMVxgz5vHwrzzyN9EfRNn1eorB4mpVFLzlU+Y8SAi6KoZDDSteDrzFXpRD7o7tAk9hDjOu2h/zZWM2CbMaanSejRZiENy3oW0KOqhHHsrTrH0lGPR/RlX5KfOp5erwelFDqdDtrtNra3t8uuoS4JjQt4oy7AcUPaqi6JkilBEbQ3Q3sps7OzmJmZwalTp0pIixIQ0Y39QTk9rl+50nPQImw4nK47D3WvPdT5AxwJY3Z2FhcuXMDRo0exuLiIPM9x7do1XL16FVevXsXt27eHAo9PDQ8p7ZN2QqPoyJRsqdomCwyCDM+dO4enn34a8/PzWFtbG/IX6vV66Ha7JQGGPp86ivhuh6jAoxli3OgsWwArR9sH/qjf61/btt3vyfL851WeH44bjfnQA4s6EeoSgR0yTajtVqewPi6AVxVoVaK7VAyFyc8nquzGyPJ+O52wMB2d0GzOwDamSeiR5yCmAXSsMboKT90Nu2XcwLnqMfyKn7B/mklQp9DtdsvqezAY3GMH/SBUzXGPMYpNR5RUP+DRzXn79m00Go0yAZ08eRJ3794tKcEh6YLgNp/a7A/hqboMu0rfWKzqpvZxcH93gxYL+/0+oijCqVOncODAAbTb7XKu9dprr2Fzc7Pcr6ElRT+ohfO1cdTgUefZ7+5o5uQb39GwW0pZnleS4pmZmUGv1yuhwxs3bpTvla6zB1mCrkpFj+q42V3JALy7EM//ci/rXuog/4V0MHheR9FiFEU81DIMUYXQjNCfz45jz41LSFV7gr4Vig/Z7ga6301smcQHa5JEZ63NhYjWGeNTOO4RpyEFYNtao3dTtfrVz/06KYYGZ35n4Hc8VN35AZUq5DoCxbgWPFzODG+IOugxTNQ+gYHUAjjnePvtt8uZxf79+/HpT38av/EbvzE0/yIKt4/dU9KhvYtQJ4w6Iz+g+HBe1fv3oVXq2OjxaQH1zJkzmJ2dhbUWN2/exJ/8yZ/g6tWrJQRKAZ2CCSVFmgXRXGDSpBN2yaFDLyVJf8ZFz3Po0CEcOXIEWmtsb2+XBcv29jYuXbqEy5cvY3l5GVEUlUKxPm04ZGztij7+Id6pS9nG6qHm/q+IfvcXehj8XJ7n3wtjDmkpZ6gj8pMQkVuyLLtHfNd/7+EMdJKgH9pz+CQG+px8+Nlfgn5Ye0PjishRRXVNnEgZ45tgLJ8moUd43O0smxbiLWNsXge7Vcm51AWdkKFWdcFVtcp0ExG8QwN/gu22trbKCzzLMjSbzTKY19kY1yWeUOwznHuNorn654Fwb5IkooAXx3GpCPH222/jU5/6FJ5++mksLi7i7t27Q4NgX48rXO71DcJC80CqNinwEH05rPb9LyJAUCdEENzTTz+NOI6xvb2N5eVlvP7667h06VL5XvyKmV4P7T75NhfjuuVxxYG/ee/vO1HgUkrh6NGj+NSnPgUpJbrd7hAkKoTAm2++ia2trXJ26IvQVlXxVQreo+JekYk+tFx0p7/aOTa78PU4bfz3vazz5a5W/ztofTaKon30eRB8S0WDv3pAiT78zKp2/MKOqWqGRI9PJBL/2gxJMnXoym5UEOriyDjFl3HXoLUWMLYDi+2ry3en7LhH3guBbRitsjrYqu6DrJL5qGKmhRdaOFz3iQn0p78AmWUZGo0GBoMB0jQtoSsKhqEIaNWFFiacMBGNw8XDPQxKnL61wWAwKIfpjUajZMRtbGwgiiJ85jOfwRe/+EV0Op17gjkFX0oq/qKmrxgQ3uihJ1NY9YVq3VShzszM4Pz58zh//jystdjc3MTly5fx7rvv4saNG0PGe77pXBXlN3QnHQeNVAV9PwH58JL//g8dOoRv+ZZvwfHjx7G5uVkmnu3tbaRpisuXL5eB1y8K6mi893m3fKDsuIlmRdtLBsDNw439/4YNtq93kP1CnuffDGDRT9i0DkFMTrpGafWBZkj+vMYnLvgdKiV7/zxS4Rh22v794TMT62DwhwGt38/PgzigjTErANvAE3w8sUmIc96xxg7CoDFqU7rOuniUGKI/0KzqlqqqMgryRD8m2Ry6kVqtVtkRhc8XKvrWVWP3M9/yu0G/K+l2uyVkRQSLy5cv4/Dhwzhy5Ajm5+fR6XSQJEnZSfhEDd9QkLohShz+e6Bz4Q+mfUiTXh9Rt/2Ee+zYMRw+fBgXLlzA4uIiXn75Zbz//vu4desWVldXy9dCr89XYKgyZfM/y7oqc5y6M31GJMtD75/YbbOzszh16hROnDiB1dXVkrZN5+jixYv40z/9U6RpOgRF+arsVfthoyrjit0VW9B4H4tlxtuD1Y0j7YWXRbfz97fR+zsqz79bRtERzjn3ZZz8HTtaAaD7gjy+fGiXChC/gPOJKD6hxb+nfYjOVx4hkVO/o6ojJ+w2EdUVyXU7Q7VfxmQMuMO52J4moQ8jCTGeMotBVXVS51EzzgBsNyybuv/22Vh+kKIbzHd5rLIL9wekdTDcpNBRFRxR1SVRUCSsPM9zXL9+HVtbW6UFQq/Xw9raWgkZ+YNbH9MnmI6ChE95JRKHT1QIt9kJlqFDKYVTp07h5MmTWFxcRBRFuHz5Ml599VWsra0NefWERoWj4JJJmXB1atkEsVJQ80VuqTtqt9s4depUyfbq9/slpJTnOd58882ScUh7VeG87mFMIRibXOLqURy3ukv9wzOLr6PL/58d2+moPP8hGUXHOOfCJ/yEdGnqOGdnZ8t5kU+Q8WHMUEl71FJ6iBjULQOPig8fhIJCeM35VPbiNwaSi+uC88E0CX0YcBxjubU2q6osfHFEvzOqg+PGdUVVQ8M6uM+HZkLNLIK+fGjBT0R1FOxRmlKjboRxA1ufTt3r9cohPwB0Oh1cv34dzz77LM6cOYM7d+5gZWVlaL8oVK6ukuj34TmfTefvMlUttWZZhlarhYMHD+K5557DoUOHoJTCnTt38PLLL+PKlStDbDwK3mEnXHVudovhh5877ZYQG44SM8FEvV4PJ0+exIkTJ3Do0CHcvn27ZErSrtWdO3dKtYSQsDFqY/5+YhljXDH2eGmL3e7czY/MHnpH9MX/Z1ttbed5/leiKDrKORchguHD3/RFquR0Psm40ZeC8jsfP6n457fOG6uu65ykYNlNN1SFdEzy82Latx2J6AoXYpqEPpQkxFnOwDJjjBFC8JCI4MNaVbORqoBUB9uMS0bh98Ivei2c83KXyNdw87uDKnilDpbzE9w4za1Rm/dSylKBgKpvYwzeeustHD9+HAsLCzh9+jTW19fLmVEVE67K+ZWWWGl+Qq/XhzmoivVnR1EU4fDhw3jxxRexb98+pGmKpaUlfPnLX8aNGzfKwO8HpjBYjZPjnwTK9Pd/KAFR0pybmyuTqE9GOXnyJD796U/j4MGD6HQ65QyQXuPS0hK+/vWvl52kb3pHzLBJlNgnT0LI8BjKutzavqMOzx6+jAH7J9v5plF5/pdlFJ30E5GfEOiaofPprwYQxExkA4LziCxSFQ/GFZ+h0d0k18/DdlSug+KNMdZqvRZFyRXOeW+ahD6cVkgxhgyAIZn6OjHJkM5ZlTzqlldHBa9JIB8f36Z5ULfbLW0hyGzOh6CqElD4nupmVnU317jOSQhRbu5ThXnz5k28//772LNnD06dOgVjDL74xS+W1TvNbXxFg6ob3F94JfjOT0K+hhgREGj+Mzc3h263iy9/+ctYWlrCxYsXsX///qHkU7WMeD+QSZ3lOwUkKh5IgcHfuid24JEjR/DSSy/hyJEjAFBaYQwGA2xtbeH27du4ePEibty4Uaol+DBlVcX+QPMHYy2AlOHxFLi8vX1bH5k7coVz8U+30o00y/P/jZTiOOciqupK/MLOV7EnMhDdVwR9+xJNxNKsgt9GiadW2YpUJa/ddE2jOh3//fpQdjAPGnBr3xOM33x/+ZadJqEPB47TALLwkw+TSd0spUpzymfbVA0JRwW1UcNueg4aXtNro4qa5kQ+jFBlNTyOoFCFc9e99/C/qYonN1ZKSpcvX8bRo0dx8OBBHDt2rKSgE7xEEFRVh+iTIXw3S//3/a15IQT279+PEydOlBpwvV4PX//61/Hqq6+i2+1i7969ZdUbWmb4CSgMNvcbGPzZFNl1JEmCZrNZdoP0e61WC9/5nd+JhYWF0h+IiB7WWly8eBEXL17E+vp66UMVirjWVeoTuqhWfeaGgQ3AHl+p/1tbt/SRuSNX5tj8P98abHQzpf+W4PaUkDKpgphp+dvfUSM3Ydono4RE3RH9jq8ZV3WfhuocoaLCKEhtN4kovMbqGLBhEirjkTE9ycRrgot1POHHk0zRNgwsx4QVXqgrFypqV9E1J3nMSQ+f7eNDhnmeD+m6hY6Qob6cTz32E2RopRCKO45KqL6Ssa9/FkURbt68iTt37uDAgQPYu3cvTp48iatXr5bkgyqXz3CZ0IewKImFMkYAsG/fPpw9exZHjx5Fu91Gv9/HpUuXcOnSpbJj8PeO/MQbzlF2k3zG/TcFNUpA1AWRAgUl1nPnzpUJiM4fQXXXrl3DG2+8UZITqAihSt5XCfA/57Dq3j3cYzVjvMcYHus9kltbt/SRPUff3cP2/lqnv7XVN9nfZUY/LYRshdczFQVUMNJumt9R0qzVZ2vS44TLryGTLnSErVOtuN9OKLxfqlyLqwqhISNAozclT14Xgvef9CTEn9gkxJnmgmcATCjYGX7A/uazT+2sG0TuwlBqZIAIKxsffqJgRkwp+vJVFvy9Gf91j+rwRkn8Vy3h+QcFw35/57rO8xx37tzB6uoqAODw4cNDqhE+m6uKlRZi6r4+F8FzeZ6j1Wrh9OnTOHLkCGZmZgAAS0tLePPNN0slgVarNTQf8DuIcE9kUpfOKjn+sAIl2wmCKomqHpJPzp8/j36/jzRNh2wc4jjGV77ylVL41WcCUlU+jsFXt+806jMuDs0YengCpP5vbd60y/2V6zPNPb/TRPzfK6Vf0yrfrus4KGH4S8O0kwegdA5uNptlF0TsRX+p2pcLog4qvKbGFSyhmkndV12CmQSm8wpMbbW5Lpi49N7q7d6D75FNO6H7heMUZzy3Izoh/8KocukMtcOqmDN1s446OG7cDKLK+4duDl9/LPQNqtrWDquwcay9uovbv9l8iIm6juvXr2NxcRH79u3DhQsXcPHiRWxvbw+Z9VXJCNHfybqBEl14U1ECOnHiBPbu3Yter4eVlRW89tprWF9fR7/fR7PZLJNQVSKuEkKd5MasOnd+IKGgJYRAs9kcSnSUnA4dOoQzZ85gz549WF5eLu0yKHGtrq5ibW2tVEnw5ZPuqXBrtvIn7eTCmZaxVoOx3pMkcLncX76x0Dz473l/e6uvB/+VteoTQsq9oZWDr/nmz10JUSB421fmoM/FZ9L5yYO6IFrIDuWyqtROws9tVMwYVQSG6EdYOHtdUJdb9hoX4jY+AseTS0xwdraKPudxN22V8RgFk7DCqvLuqbvh63D8qucPkxzdIACwvb1dDlV9yfsqGNG/iMPk6icv/9+FiaEuUdH7oapda421tTVcvXoVe/fuxQsvvIBz587hj//4jyvPWUg391lLfufnO6GeOHECL774ImZnZ7G1tYWrV6/izTffxNLSUskc8xXLwwXEus96EmiuCu70LQZIzZrkgOh3aPB9+PBhvPDCC/9/9r4kNq4sy+68P8QcDA5SkBQpZpaUopQjkFmoAlxVgNMF25veGl41YAMNNAyjAbt7bcCrWndvvPEIGL0x0AaqXQa6AVfDKFRnpjM7s9SZpUyxVKRKosQpOEaQET/iD+95Qd6XL77+FMGgpKDeBQiJwRj/j//Ou+eeey7eeusttFotCbIE5q1WC59//vkzt6vihkG+u2m3PXO7EAE7BaGxsnVpOLuNerH+qdWzfnLMT/5t4Hn/wLTtq+HNTrinR128aRNAQphisYhcLieBiP5Vvy8EYHGO3eprpW1C4+rDcQMswxlTlCABAALPPyyY1t9ZptnSIPSCi0KMMR7OhJLGI4TVNeEvVNSXI4HmiLxvlkJkONui+ThU96A6gkojxlkMpal60ixoohyFqSt9YmJCgtzm5iZs28by8jKWlpawtraGo6MjCSiUxalFX/LnUjl2WhxKpRKmpqawuLiIN954A6VSSbpgP3z4EPv7+zBNEycnJ/L4qOcwzt8vzcw16nyEi8AERI7jwDAMeRzoeai+tbi4iA8//BAzMzOyV4VqWY7jYH9/H19//TVWV1elkEOdRRV29Y6jVaJMONNoReV3n8FwGMPYWf03nMb+fGXuC6Nr/KTlt/7Ic91/Yudyc3HqxbC3nvp9VqXcJCohii6KRlZrQYNY9CTViKJERmkgFJEteQiCR/lC6esnRw1Hg9CLxaDTf5A+oz6OogsvwMPQOAPQh8/0IKh1EpI7qz5zqptCFAipA/iivtyDuEGEwVjNyoQQaLfb2Nvbg+d5WFxcxM2bN/H111/L4roKMGEqk+5DgOY4DmZnZ3Hjxg0sLS3JRfzLL7/EgwcPpJmn67rodDq4cuUKisWi5PLVZtmkabhZACi8MKjUKGMM1WpV9iSpnnv1eh0//vGPZY2s2WyiUCjImtC9e/fQaDTw5MkTmb3RhFqaapuYwQwRMc8RgLEuxnT889bJdmu+Ov816xp/2vKOjn3X/T3DspYMw2BJG8I4qkylkCkbV9sH1JpiuMUjbZMbZk2yZLep1jzh5+H82DbMv7Ut6ykuSYytMOEsE2JxxdtwL0EWcEpzuB1ErJBGlYS5Y6KayOKHqIKonXDaKPAshdSoTEg9hlQPUW1mTNNEq9XC5OQkJiYmIrOxsPBDpdJM05R9NvV6HdeuXUOtVoMQQtJwNAhQ5eZpoVCztbh6W9aNSNR4DFLxUVan0oe0aAkhUC6XpZO3EAKdTqdvSNvu7q4cqqeOkCY/wSgAytoMOUQEjDGPjSkIAcDW8Va7WCx+U8tN/gcT+K+B768Kwf2486lmEkSdhqfzRqkPo/5Va4RJatg4Gi3LOjMICHHf383b+U9My2peFhAa45oQ2BmIsigASqrLxPG54awiKesZ1M49TpEXdj4ghRothOE5KoPMHYoDorTdHAF3t9uVIEB2NI8fP0a9Xu8DoSgqhG7vdDpynDhx9N/5zndw584dTE9PQwgBx3Hw6aefSuduWiA8z0O5XJZ0H/WGhEEubZeaBEDqqAA1AyL1YnjYWj6fx61bt/D+++/LzJCe13EceJ6HX/3qV2i1WgiCQDqTk0qOakqqQCNrxpaUkccOcRTgjDEfDGPd0LjR2uotTMyvQODPO97JvuP5f2iZ5huGaZbC32s1u4mq86qb1LhrYJBa3KDZ6TDgAwA8CDpMiC8tI/fg0f52V4PQSxACYOrIriggilOQRV34akE/jsqKm7g6rIw7PGaB6Bo1G1IH4YXfU9TArUF46ziQpqyF7mfbNprNJu7evYubN2+iXq/j+vXr2NzcRLPZ7DMtDc8XosW81+vh9ddfx3vvvYd6vS4bOakXSZ2qSWMNJiYm+qz3VUfjOEFIeKcZNRYhyteOKMh8Po9KpdLXj+S6LqampvDmm2/iu9/9bt9IavIC7PV6+PnPf47t7W25yNF4b9d1pYVM1A48SaBwPqpO+AwsYGBi3BerjdYWB/CwXpj+KbqtQyfw/9iEuG2aVjV8zYdVn+Em1DhvwbAoKaqWk7TxTFKopoFQUqYOACIIdnOG/TeWZe3gEsU4g5AhhDCNU6/6yHkxYaoozjUhjs9VC5PDNKXF7YCS5NK0k1NVYGotIiwrVWta6vOp81aiLpIwGIV7kOjzdzodlEol5PN5HB0dYWdnB6urq3j33XexvLwM13XlKIUoubdaGH7nnXfw7rvv4vr163Ig3ebmJu7du9cn4aYsSK2dqKM0ogrGcYq/sGdYWIquupsLIWRfiSrzdRwHU1NTuH37Nt5++23ZtU/AS8d7a2sLW1tb8nwEQSDdEqh5NdxbFLehSTKyjNvkRC90CAD4APhlWbQa3YONemH650b3uNUOvD8R3H3HsnNXozadYTYi7hpPum9YvJC08Yl7vjSbnig6r+89+L4D3/+qWJj49MnRTkuD0EtCxzHANBIMNMO3pWn3B50ffx4wShvxrRby6ULIKsAIe2INSx+QmzUp08jtoNVqQQghrXyePn0q5wSpj6fsgmip69evY3FxEZZlodls4smTJ1hdXe1buDnnaLfb6PV6qFarsqYSBp44n7ooKb662aCLmyhPAnmq9ZTL5b6eE845qtUqPvjgA8zPzwM49YOjnh/Kdg4PD6WzN410UC19VDHFMOflPDUhAGNPx0UAUWOufPVvzfbx0bHo/pHnuj84m0tkxg2pHAbMwxvYuJaHJFFTXA03ampyXFNr4Hu7BVh/ZVn2E1yyGF9hgoAhIKzT7wBLTI1VikkVK4R/oui8i1os0na4Km+dRaKb9BpJM+qj6Dn1GKg9MzRrqNFooNPpoFAoYGFhAbOzs320IXWu0zC/SqWCpaUlTE9Py2F+W1tbWFlZwcbGRp/1DanTut1upCN50k40LutTqbfwDwFFPp+XogFaDDzPQ6VSwZ07d7C4uIhSqSTdEAjcHMfB1tYWvvnmG6yvr8vHdrtdqQokOjKpJneBHe8BYwge722Ly7Z4bbd3j8qViS9qrPwTC/hvvufd50HQThvPHXZRGaRGM+j9k+TYcRRxRC3IYV7w93k7/8snzcbBZTuPY5wJCePs/bO4BTSOokvLhC7sHQ/IDVMWQLWHtIU3bix5Uj0rbkYSvbYqTSaA2Nrakmank5OTmJychOu6crGl7IcK8NeuXcPNmzdRqVRkjWR9fR1Pnz6VDsjqZyG5ehwIDXKuyCKIjqEqw6YMKJfLSQBSj0epVML169dx48YN5HI52fNUqVTkuPONjQ08fPhQNtZSZkSLiTr1My4DvlC6AAgAFuCSxtZJw1mszX9tdexWxzv5bdf3/7UQ/I5hWlNRlGd4MGFcHTk8giWcaWdtCUnacIb94uKcUETgb9uG+Zd2LvcE3ct3DscWhERIHRdVIwiDUFyHfZYv0KgAKlMBMsLPLG73HLWzSqqBZaUSwxNPKVs0TRPNZhOPHj3C9PQ0GGMoFotysVcLu5xzXLlyBbdv38bNmzel7c3u7i729/efoRzV/iQabxHnkZZWd4uiT1QAIvl5oVCQdSDV2dw0TVy9elU6OTSbTQlMjuOgVCrh/v37WFlZwe7urjTPDDuLh7311M1BlKDkAgAqOAWiyxtPm1scwON6ftqxes52O3D+jRe437Vzufk0hiBuBErcpi6K+s068iXp37h1gAf+sRHwz8qF6icbrb3mZTx/40zHQQhhgCVnNHFZUNzwuTAtF3Vb1PMMC0ZZRzQMMiMnjQpIy9DULIJ2g2S4CQC9Xg8rKys4OjqCEAKzs7NYWFiQu0u1tmNZFmq1Gmq1GnK5HDY3N/HJJ5/g4OBAquBU4FQbUpOy26zHVDW47PV6fZLxSqWCiYkJFAoF6e7gui6q1Spu3LiBH/zgB8jn87IRtVAoSMXgwcEBfv3rX2NnZ0e+Fj2ehAqkhksyuL3gzFuc1YQuNQjJOlHvoFEuVz+bMCr/ngH/y3Xd9ah+oj6qK2JuTxxdF/f/YX7CpsqxrQOuu5G38v8zl889vaznbZzpuDO2YXAESLN2SVvo4upPabLMtJ2ReqGEueGoeUVRjbhxdZM0c8XwMD9V7UNUluqrdXJygna7jcnJSczNzeH111/H7u6ufKznebAsC1NTU5icnJTmkSsrK1hbW5PUHdnhUBZEBXySR4clzYOAu+qCrQKEbdsol8vSt4+yI845ZmZm8Oabb+LWrVuwbRudTucZQ9J2u41f/OIX2NzclO+VQE615KEsKG3zcMFgxF8VEAKArXajNV+ZvSfa+LO2OFnzPP/3TSN4zbJztaTWhLC6Tc1W0wZjRtHZWdmPJDDzPXfXDMRfF4rF/7d+2DjWIPQSRN+FCxgCMNOyhHBWE7VQD2LXk3UhHNQFOUkxl1S8zpolDHqcVck2yaVVsOWc48mTJ7BtG9evX0elUpE9PvSe6/U67ty5g2q1Kr3U9vf35cVN9BWp0brdLvL5vGyQPS/lSQKBcBNqoVCQIKguPpVKBbdu3cKtW7eQz+flaG6VXjs8PMRnn32Gzc1NFAoFeJ4Hx3H61IuWZcler/AmZRRS/wF3agG7RPLsTEB0suMCWJnJTbY6bvt3Dvf+Fe/13rZsey6uJSNt8xh1TQ9SD0raaEZmQUHQYX5wt1Ko/IVlW9vjPKrhEtNxwjAYs4QQRtrU06QvRHg0dBz9lrTYx/2ehToKT4ENp+nh3Zn6GuquLI4yzPJe0ujKcHHftm24rou1tTXs7Jz2zZG8WaXXarUarly5IsUK6+vraDabfY7S9Pnz+Twcx5EZySDHPUpkQRSi6opN9R/qP6LXpixnYWEBy8vLcqqsekyPj4/lYLqtra2+c+e6rrQjKhQK0hkh3DMSJ/dNq0kMs8GQoHcGRHgFY9892qwUJv5PBYV/B+AvPc/7reBBO4meS1KrJf2elZ5LG4QpWzI8dz3P7D/P2flv1g92vMt8nsZZmGAKRR03LA0XRafFNbGGQSOJXknqS0rqUUjaIUcBTNzznycrinp9kjhT1uK6Lo6OjtBsNqWQoF6vo91uy8WfxoQDp7Wex48f4/DwEJVK5RnFEdF3akNnmhNE1CCxKOt9UrSpFCCp92h+E+ccc3NzmJ6elu7guVxOTpnd2dnBysoKDg4OpFqQZNgkZKCxAc+xByhLJvRK0XHh2O3uN+cq9S9Mx9rtBc7nXT/4l4YfvGHn87NZ6dBwo3NUZjPIOY/KhFQA8nq9HYuzvy6Xy7982to9vOznaHxrQkKYgLDYgFd8UkNr0v+H2YXGKWiidrtZQSFr/1KaNc+gFw75uRUKBbmwdzodNJtNNJtNVCoVLC4uYn19XVr1LCwsoF6vw3EcnJycyB4bkixTHw0AtNttScUlmZQ+k8qfAVZYeUZAKYSQ4gPVhofAiGTaH3zwAd544w3s7+9LUCVfuLW1Ndy7d0/WvMjVgUZvEPgQgKoL13lp3bSsKQsdh1eMjgvH9knDA7A2k5ts2q5zv4Pev+j1ev/YssyrpmlV0ijyKEo/nK0nXctRNWDVhaG/DuS1mB98VilW/8Kyrc1X4fyMcSYkTMaYlZVbTwKdLKOw47KmqN1Q1EKfZDGTBBxpdvBZFGNZQCdJcEHZT1iqDQCtVgvb29t4++23Zb+QEALXrl3DzMwMDMNAu93G4eGh3P0RdUWgQPUgypBU1+ysPnhh6o6ynEKhgHK53E9RnWVe3W4X09PT+P73v4/l5WW026dMTS6XQ7vdltZC9+/fx87OjhwpTvOCAEhADQPQMJuWuM81fD3gTB03xg7aI6bn9ubKV1tW19noBO2Pe37wB9wP3rByuasAzEGuzziqPrz5iOr9iVXDBUGXe979aq70nwr5wpfrhw1Xg9DLjUJExw18wSeBTxztlXUhCC/6UW7cUTunLK7Pcbu00SWX6TQg1UnUDISyokKhgJs3b2J1dVU2gZKwgax4fN+XjZ/UpEqvQcAWR0tGNQuqvUlhw0rDMFAulyWlFqYU5+bm8MMf/hALCwtStk3HulqtYm9vDx999JEcyRC2QyJXb3UA2qCAEaWqPGf207dTE4DPXmE67pmsqL3rAnh0JTf5U8ttr/Tg/TPPdf+pwXDNtHMzcecwPFo8qRk+bUMRNS1VcN4N3N5vCsz6z8V88ZP1o8bJq3JOxjcTEsIcxfvPmh1lXbjDABTnYRdH2w0DGMPKfbN46SV5tHHOcXBwgEajgeXlZVSrVczOzmJjYwOVSkXWWo6Pj/G73/0OzWazj9ojRwVSrUUN8UvaVSbVgCgTImAiqTY5IywtLeGtt97ClStX+sQQ5Hi9ubmJx48fy6ZakmuTeIIGEaoTV+NqiufZEMSJGjJ+PwUumXnpqGLPPTqaK1/5u7zrPel5nb/pCu+fu677I9Mw6qZlTcRtENQ6ZXhCcpbzGa4DAUDg+13uug+KRu4/VoqVn20e7++9SudinEHIhsHs5/A6Ay3QcZlQ3GiJKCCJ+z1q8R3EBWKYelDUIq/WbNrtNnZ2duTU0MnJSQko6rRYIYRUyu3t7cmMiFSAJMtWsxGyunnGxiRk9BqVKVK20+v15DhniqmpKXzve9/DwsKCNDD1fR/FYhG9Xg+NRgONRgNra2t9Kjt6Dtu2USqVzpUxZ73/OW1+CIR0RGZFewGAjdnSzEGu13vQDZwPujz4/cB13zEYaqZl1QzDtOLGiEdtKrOMFglRcE3uur8pMOu/VArln22eHOy8audhfEGIcxvGxb3/YUd8x2VCWXfJtHhGfanj6h9pCrzzUnYqxUV0luqFRqMPaHGenp5GpVJBoVCA67pYXFzE/Py8BKSPP/4Ya2trUmXmeZ7MiFQbnzDHHjfePHx8LcuSRqmkXqPenW63i5mZGSwtLcFxHHQ6HdlY2ul0cHx8jAcPHuDhw4dSQk41Iqp3kXgi7ti+LD0djDFxRsUJ6IiNnc6+A2CtXpxuFFz3y17QfccV/j8KPP/7nPnzhmlNMcOopG3skqi8MN3Kg8DlvrdjCnxesgr/vVQsfbRxfLD7Kh7/cXZMKAKwaYEJp8RxM4XiFtms5qZxKreoHpC4jCLcm6TONokaO6zWIVRASAKhrKOu08BVXfhJskzjt0ulEm7fvo0PP/wQpmmiWq1ibm4O7733nmwUBYDZ2VmpTnv06BHefPNNtNtt7O6eXnOO46BcLsusQxUXZDnu6sCyqOmwav8SCQsODw9Rq9Wk1xtjDJ1OB3fv3sXa2pqs+QRBIJV9pmlKTzsC46TJmWk0aVjAkNYzFJd5R4kY5DEBOF4eyfhLHQ3n4BjA8dXC9NO8733q++53POG95/n+PxTAMmOYATMmDMMoGaZpR2WqqdebEA73/QPueQ9smP+7mCv8Ip8v/HbjeL/1qh738QUhhgpjw9NxgzQBZqFcsowAT3tMUqaTBGqjyHayHCtSyOVyOUxNTeHdd9/FjRs3MD8/j/n5eRweHuLg4ACu6/b1C6nO3JQxqaCa1CB8HrqUlGutVguTk5PyMzQaDWxsbKBYLEpPvIODA9y9exePHz+Wmxqi8wh4SZpN9j1j0sUudBo0WOx2DzoAOvOVK1u+7//a9/2/8gP/tZ7o3uGCvx9wvhz4/hxjqBqmWWaGkWfMsA3DsCJECT4EdwXnbXC+j0A8yJnWR/l8+aOcnfuNZVsH64e7r3TNbixBaL42Z3Y6zSoYy2V1gx50wc5SsE97XBb12yjAYVBabdhBd2qBXwiBWq2GfD6Pzc1NPHnypO91SDl2fHws+20A9NVSVI+1KCv98wYJCqgmRc99cnKC1dVVVCoVCCGwu7uLjY0NPH78WNanHMeRTgqGYSCXy0mboYs+r6MEIGg6bujYOtnjAJoAmrOVmUd5v/CF4P7PeBBc5SKY9bl3y/eD2xzBYgBMMaAAIIdTJxoBwAXQNoFtmxkrOdP+yspZq5ad2zRts/XkaE/X68YVhITgOc75rGGcbk2jxnsPstiO0nMtSpIdR8clecHFgcwoM56sz0V1Gvoh5RndTpQW/Z382UiC3Ww2EQSBlGyT6ICUZZRhZLVfisuEotSItm1LS6BSqQTTNOH7PhqNBr766isAp71OR0dHErTICYEyHrWBVp2zNAZXCqDl2SOJnZN9AeD47GdjYWLGCoLg48APCkEQlHnAS1zwIoA8wEwGCMbQMw2jY1nmsWXbx5Zldh4f7fXgtvUBHXsQ4twWQtTDdFyS28EgWUPWTCktG8oiv85Si4qaRzPM+xo2VEcCtRdHpeiofkMUVqFQQKlU6nOSJmqu3W73SagJhMLgMqxMPmpMOhmZkq+b4zhyEirZ+NBAOhIz0HuzLEv2Q5GCL1y7e1kvFQZ4OhMafWy09n0FlHYT89AAQE8fs0sGQsISENOGYVg4J7U2ikwiSYwwbB+QuqBGybrTxpmP8hio9RvKduj/qv1NuHGTRnST9JkW+PX1dTQaDUnNxVncDLJpiDsHZI5KwEMmo2qtiuyDPM9Dp9PpsxaiURLhcedjcZ1IEGIahHRoEBrpzlxwG0CNMWYJpNdvRk1PDZp9xHXEx1FQg7zuMO7Kg35Wdcy4OhKZ/m9Zliz8U6Hf9320221wznF0dISDgwNsbm6i3W5ja2sLlmXJ+ybVg7Ien6RzQJQa0WxksaPen2x86L2QxFtV3qkZ6XMaxXDuS4WBuWC6WVWHBqHR7vCEyAmGKjMMS4R2pqO2shnhex5ocX2ZFjg1a6AMwXVdbGxsSOFBu93G66+/juvXr/dlSADw9OlTfPHFF1JZR6O0AfRZ4UfJj4c91sC3jbzU31Mul+G6Lk5OTuR7IDqx3W7DMAzUarVnMj71/BEQqfLxlzgV4oyxLoP2jtOhQWjUC3rRMI2KEMKMssUJ98jEiRbimkGzOGmf1yMsPDguLlMaJKNKGlER5eSQJHpQ70O3hymslZUVKUwAgKOjI9TrddRqNVkzMQwDS0tL0saHnBS2trbw6NEj7OzsSDosLCzIUhdKclFQHbNV0KMpqwRQJJooFAryWEbNAsrSD5I2MG3Um4s4J47TfzmHYA60OEGHBqGRg1BBgBVGQaUlUXIXpZp7HjHKjJAWT7VAL4RAp9ORdaCJiQlMTEz0jecmKXe1WpVO1lTcr9Vq0iRUlXAPm/Wk3RZW5akgSS7Yg44SH4PgjDFHu2jr0CA0ehDKCybsLIvtIAalw9SPXgbaLKtq7rwgGqaiTNPE/Pw8lpeXMTk5iXK5jGq1+oy1PanMVIudXC4nJdxZxlUM+reo909Zci6Xk8BHt5GKT6UGx6Tuk0THBYyxHtPqOB0ahEYPQkwxL00bZx1XjB+FmiwrGIWVbarK6rzO18+jYZV6giiDUF0TfvSjH+Hw8LDPHZvoLsuysL29jadPn2Jqagqzs7OSvgs7Eg8LlGmzX9RJlqqTQph2Uym8F1XvGTFlJxiYB+2irUOD0Ki5JhTATt97kv3OsM4IaaO7s4DRRe2i1R36qPue4oAzyhHcMAzU63WUy2Vsb2+j2+3KqatEeVGsrq7io48+wu3btzE9PY1cLodSqYRSqdSnUksaTxEnWshiGBmXBYc/V9xAsjEODsAD0xJtHRqERhbzU9eY0z4uGoZhxXmNJWVBWY1K0wAqbcRD1r8NkwGMytYma2YXBh/KGKioD5wW+EulEvL5PFzXheM4aLfbcBwHx8fHmJmZwcLCAmq1GjqdjlSfpYkwhrUYCh8rlR5UgTVuTPNFA1DYkDTsCD6a1xeCMeZrOk6HBqHRXr22gKgCzB52lz+ONaEotVpcVjTo50j7DKpDADV1+r6PnZ0dORYBgJRgG4YB13Vx//59dLtdTE1NoVAoYGlpCVNTU309OcMAb1YDWZkOhFRySX0+Lzr7GfHrc5zOE9IgpEOD0AivUgvAFBjsrIAzTNYzTLf+sIv8oIsTqbyed91C/Sy+7+Pk5KQPTNSJprZt49q1a2CMYXJyEq7r4rXXXsPk5CT29vb6mkAvYiGPGjoWR/eFe5YuhSgBAAQEA9MGpjo0CI12geEmIKYAmOqEwrghb2mz4IcxPM1CGyX15cTRMOHsJqq2EberjwKM8GIaN4AtqQ5CDZ2qe4BhGPB9X9rh0P0oQyLRwszMjHy8bdtysJ3neX39XFHHa9AsIa2elOTnF+c9F3efqFlL6jmLO6ZJI7rPOwo85vGCMXDGNAjp0CA0yl2uxQWvgpnWIJnOoJTdKOmsUWch4eF9wzzXsO9BXTBJLUfgQ42rNCWVbiPw2tvbQ7fblXY+cZnoRWRI4yKlH+Z8JHwHBXQmpEOD0MgzIeNsoJ0Rzn4GqYsMWzeJqktEUT7hXX1c7WbYxVbNIrJSU+c9DupnJnCh+g6p4ciklNwRhBByNo/qP5fP56Vb9UUt8lmcJ14EAF3U60eAkWAAh9AgpEOD0CivZgtAhTFmZV3Mh6Xbhh1sl3afi8yeLir7U8E1TGFSoyc5ZXPO4TiOBCYSNVCjKwFo2Lw07vXGHYCiXv+isqKI4DoT0qFBaITBeWALiAozDPMiX+c8fUcXtdCMCjxHtZjS2AaywVFdCIBvRyRQ5qSCWJI8+3lkI5clUj6TOP3RE751vLxhjNsbDoIgD4jKsAB63npI0t/PI3AY5v08LxVXWEAQXgBVx2y6nUCHFHNht4iwYGCUC7HQa27oeOhjoENnQqO7oDgvCgMVxtjQmdCo6kXPU5QQ7hM67wJ+nl6iKDdp9bbwELw4UcXzzG4uKzCl9KsxIcA0KOvQmdBoowyGYtwCGLVbD0tqw6KC88yxOY+PW9bO+LgFPur382Z8WT6r+tyu68J13T4Jd/g4Rn1OovDCjxmlbc6gnnxxvyeJCqK+g0kS86jvYNr4jnAbQtLfQt8L42yjyfRSp0OD0Oh2vhWw/jEOrwIFE6W+u4jPnZRhhQ1HiXbzfb9vhlPUQhuuDWVR9w0ysfZ5ZVQv8twPcTYNAWELIQzo0KFBaGRXZI2dgdConAjGEcBGQcmNMsKu4FESdnXHTnWky9gP9PJ8SWAIAQtCZ0I6NAiNJOaK05ZgmGOM5S4afF62xSyqE3/UGVFS82jc/ZMymqiMiB5nmiZyuVwmFeKwHm8v/fjt5xOm0HScjpc4xkuYwHlOCDHPDCP1fUeNVIizsImy03kRWU3cYhtXh3iRGVjcbWkj0tUsKGmS6XkslHTQAYEA0x7aOnQmNMpswIYQNQDGMFRUWvE3fJ+XeVEbNRAlZSRhgKH+IADSAUHNiFSqkO5LwEM/WZt9o86FBpvMGNRjYA5jeqidDg1Co3qz7CyCrAtp2oI1LjWhF1n/icp81JlCvV4Ppmk+44RAwBMFQBpMLhiAOO8ygYbJ2N5O+9DTR0SHBqERhGkYvmWYmwj4EQ+CE6GsYqPKioa93wVlfqmAMIraVprDQtzfySWBxjmoCjkAEoCiLH/iXMcH3TDouk8kADk8CBo2rLs5y97UR0THyxxjVRN62j08mbNr/9cLghsc/H0hUOcCOWaZFgzD5N9mSjAMQ4AxMINB8FN63DAMSY+fLYSMMQYBuSiy0z8xADAM4/TXs4WPPcN2xCz2QnAQQApx6h4ZBAEE/1bWrLhLCyGE4DwQUvYccMY5Bw8CdnY/EQQ+hIAwTRPMNEXgecI0TQEAXAihrsXG2Thn+kycK44HZ59PAGAGe/aDhDCIPrfggl6B+b4HCMCwbc59j4vAF6ZhFG3LFBBcGIbBuBAGY2CcB9wyDWEYBj89qMwwDJNZBvMZDzoi8E3ueQYTgjEhGDMYwBhOR1KzzH1UMe899cGccxZ+njO/z2dvF6fHQPk+iNPb1MxO7RcyzoCT03kXZ98BoYyUEPz0PoJzDsGFUOXvZ0999rrfvgf2zCEQnHPhC847TKBRZLm/z9n2T/M5exM9vdDpeIlZnh/+j18+BpDTh0KHDh06dDzncC0ACwBMfSx06NChQ8dzjsAA0NbHQYcOHTp0vIBoazsPHTp06NDxwkKDkA4dOnTo0CCkQ4cOHTo0COnQoUOHDh0ahHTo0KFDx6sBQmV9GHTo0KFDxwuIsgVgA7pZVYcOHTp0PP9w//8ATHPqr1bJ+qAAAAAASUVORK5CYII="/>
</defs>
</svg>